MZP      ��  �       @    �pjr                             � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                                                                                                                                                                                                                                                                                        PE  L ��b        � #                        @                      `                                                     @                                                                                                         .text                                `.data                            @  �.rsrc    @      @                @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �pVT          @  �   `  �   �  �
   � �    �   0 �    �pVT          H �   ` �    �pVT       y  x �y  � �y  � �    �pVT      �    � �   � �   � �    �	     �
   8 �   P �   h �   � �   � �   � �   � �   � �   � �   	 �   (	 �   @	 �   X	 �   p	 �   �	 �   �	 �   �	 �   �	 �   �	 �    
 �    
 �!   0
 �"   H
 �#   `
 �$   x
 �&   �
 �'   �
 �(   �
 �,   �
 �-   �
 �.    �/     �0   8 �E   P �F   h �G   � �H   � �I   � �J   � �K   � �L   � �R    �S   ( �T   @ �U   X �V   p �X   � �Y   � �\   � �]   � �^   � �_     �`    �a   0 �b   H �c   ` �d   x �e   � �f   � �g   � �h   � �i   � �j    �k     �l   8 �m   P �n   h �o   � �p   � �q   � �r   � �s   � �t   � �u    �w   ( �x   @ �y   X �z   p �{   � �|   � �}   � �~   � �   � ��     ��    ��   0 ��   H ��   ` ��   x ��   � ��   � ��   � �9  � �:  � �;   �<    �=  8 �>  P �x  h �y  � �z  � �  � �  � �  � �  � �   �  ( �  @ �  X ��  p ��  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � ��   ��  ( ��  @ ��  X ��  p ��  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    �   8 �    �pVT    (   �( �P ��( �h ��( �� ��( �� ��( �� �) �� �0) �� �^) �� ��) � ��) �( ��) �@ �* �X �"* �p �P* �� �p* �� ��* �� ��* �� ��* �� �+ �  �4+ � �Z+ �0 ��+ �H ��+ �` ��+ �x ��+ �� �, �� �2, �� �\, �� ��, �� ��, � ��, �  ��, �8 �- �P �,- �h �N- �� �r- �� ��- �� ��- �� ��- �� �. �� �    �pVT       y   �    �pVT          ( �    �pVT         @      �pVT         P      �pVT         `      �pVT         p      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT                �pVT               �pVT                �pVT         0      �pVT         @      �pVT         P      �pVT         `      �pVT         p      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT                �pVT               �pVT                �pVT         0      �pVT         @      �pVT         P      �pVT         `      �pVT         p      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT                �pVT               �pVT                �pVT         0      �pVT         @      �pVT         P      �pVT         `      �pVT         p      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT                �pVT               �pVT                �pVT         0      �pVT         @      �pVT         P      �pVT         `      �pVT         p      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT         �      �pVT                 �pVT                �pVT                 �pVT         0       �pVT         @       �pVT         P       �pVT         `       �pVT         p       �pVT         �       �pVT         �       �pVT         �       �pVT         �       �pVT         �       �pVT         �       �pVT         �       �pVT         �       �pVT          !      �pVT         !      �pVT          !      �pVT         0!      �pVT         @!      �pVT         P!      �pVT         `!      �pVT         p!      �pVT         �!      �pVT         �!      �pVT         �!      �pVT         �!      �pVT         �!      �pVT         �!      �pVT         �!      �pVT         �!      �pVT          "      �pVT         "      �pVT          "      �pVT         0"      �pVT         @"      �pVT         P"      �pVT         `"      �pVT         p"      �pVT         �"      �pVT         �"      �pVT         �"      �pVT         �"      �pVT         �"      �pVT         �"      �pVT         �"      �pVT         �"      �pVT          #      �pVT         #      �pVT          #      �pVT         0#      �pVT         @#      �pVT         P#      �pVT         `#      �pVT         p#      �pVT         �#      �pVT         �#      �pVT         �#      �pVT         �#      �pVT         �#      �pVT         �#      �pVT         �#      �pVT         �#      �pVT          $      �pVT         $      �pVT          $      �pVT         0$      �pVT         @$      �pVT         P$      �pVT         `$      �pVT         p$      �pVT         �$      �pVT         �$      �pVT         �$      �pVT         �$      �pVT         �$      �pVT         �$      �pVT         �$      �pVT         �$      �pVT          %      �pVT         %      �pVT          %      �pVT         0%      �pVT         @%      �pVT         P%      �pVT         `%      �pVT         p%      �pVT         �%      �pVT         �%      �pVT         �%      �pVT         �%      �pVT         �%      �pVT         �%      �pVT         �%      �pVT           �%      �pVT            &      �pVT           &      �pVT            &      �pVT           0&      �pVT           @&      �pVT           P&      �pVT           `&      �pVT           p&      �pVT           �&      �pVT           �&      �pVT           �&      �pVT           �&      �pVT           �&      �pVT           �&      �pVT           �&      �pVT           �&      �pVT            '      �pVT           '      �pVT            '      �pVT           0'      �pVT           @'      �pVT           P'      �pVT           `'      �pVT           p'      �pVT           �'      �pVT           �'      �pVT           �'      �pVT           �'      �pVT           �'      �pVT           �'      �pVT           �'      �pVT           �'      �pVT            (      �pVT           (      �pVT            (      �pVT           0(      �pVT           @(      �pVT           P(      �pVT           `(      �pVT         p(      �pVT       	  �(  HN  4          |O  �           0P  �           �P  l          TR  D          �S  %          �x  J          ��  J          ��  V          D�            d�  v          ��  �          ��  ^          <�  �          �  �          ��            ��  �          d�  j          ��  &          �            �          � v          $ �          � ~          8! 2          l$ �          ,( P          |+ &          �. �          �2 �          |5 r          �8 �          �> |          \B �          ,G �          �H �          �J �          \M �          O �          �P �          �W �          �_ R          �e f           Pf �           $g d          �j 4          �r \           :          T� f          �� &          � �          ؗ �          �� h          $� V          |� �          �           � \          t� p          ��           �� �          �� �          �� �          � \	          x� L          �� �          � �          P R          � �           � F          �            � v           H ,          t �            �          � �          h �           �          �! �          �% �          `'           l) j          �0 "          �2 N          L7 X          �9 H          �: 
          �@ �          �D �          tG �          4J �          4M �           N           (P            (R Z          �S p          �U (          X l           �X �           TY &           |Y �           HZ �          �^ �           �_ (          �c .          l p	          �u �          �} �	          X� r           ̇            ̎ "          � x           h� >           �� J          �� �          �� �          $� �           � �           �� �          p� d          Ԧ           �           � 2          @� r          �� �          x� �          L�           T� �	          0� 8	          h� �          X� �           T� F          �� �          �� n          �� �          ��           �� �          �� �          h� N
          � ,	          � H          ,           @ �          4 "          X �           ( �           � �          �           �  X          ($           8' <          t* *          �. \          �1 0          ,6 0          \< X          �@ h          D 0          LG           \K h          �O >          T �          �X �          �\ �          P_ �          c           e �           �e F          0h �          �i v          @m            @q �           u            0u �
          � �          Ԓ �          ��  R         �� -          � �          �� �
          � �          p �          0! �
          , �          �.           �M �          xZ �X         (�	 \          ��	 ��           v
 ?          `�
 �          �
 �          `�
 �          �
 ]          l�
 ج          De ��         �#           % A         T2 N          �B �          � ,+         �G `          4Z �          �` �         �o h�            v_          xe �	          $o �6         ̥ �          �� \2         �� �          �� �j          �\ "           �\ @           D V C L A L  T A B O U T D I A L O G  T A U T H E N T I C A T E F O R M  T C L E A N U P D I A L O G  T C O N S O L E D I A L O G  T C O P Y D I A L O G  T C O P Y P A R A M C U S T O M D I A L O G  T C O P Y P A R A M P R E S E T D I A L O G  T C O P Y P A R A M S F R A M E  T C R E A T E D I R E C T O R Y D I A L O G  T C U S T O M C O M M A N D D I A L O G  T C U S T O M D I A L O G  T C U S T O M S C P E X P L O R E R F O R M  T E D I T M A S K D I A L O G  T E D I T O R F O R M  T E D I T O R P R E F E R E N C E S D I A L O G  T F I L E F I N D D I A L O G  T F I L E S Y S T E M I N F O D I A L O G  T F U L L S Y N C H R O N I Z E D I A L O G  T G E N E R A T E U R L D I A L O G  T I M P O R T S E S S I O N S D I A L O G  T L I C E N S E D I A L O G  T L O C A T I O N P R O F I L E S D I A L O G  T L O G I N D I A L O G  T M E S S A G E F O R M  T N O N V I S U A L D A T A M O D U L E  T O P E N D I R E C T O R Y D I A L O G  T P R E F E R E N C E S D I A L O G  T P R O G R E S S F O R M  T P R O P E R T I E S D I A L O G  T R E M O T E T R A N S F E R D I A L O G  T R I G H T S F R A M E  T S C P C O M M A N D E R F O R M  T S C P E X P L O R E R F O R M  T S E L E C T M A S K D I A L O G  T S I T E A D V A N C E D D I A L O G  T S Y M L I N K D I A L O G  T S Y N C H R O N I Z E C H E C K L I S T D I A L O G  T S Y N C H R O N I Z E D I A L O G  T S Y N C H R O N I Z E P R O G R E S S F O R M   (       @                                ���                                  8   0   p   `   �   �  �  �  �  �  �  �  �  �  �                                 ����������������������������������������������������?��?��?� �?�  ?�  �p ���������������������������  (                �                       ��� �  �  ��  �H  �x  �H  ��  �d  ��  �)  �9  �  ��  �|  �   �   �  �  x  0�  �  �         !              �  �  ?�  (      
         P                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �����  �����  �www�  �  �  ����  �  �  �����  �����  �����          (   '                                    �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                     ����� ����  ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ����  �����                     (   !            �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �����������������   ������������wwww�   ������������w�ww�   ������� ���x�ww�   �������  ������w�   ������� ���x�w�   ��������� ���w���   ��������� ��wwx��   ������������www��   ������������wwww�   �����������������     �F o r t s � t t   a t t   a n s l u t a   t i l l   e n   o k � n d   s e r v e r   o c h   l � g g   t i l l   d e s s   v � r d n y c k e l   t i l l   e n   c a c h e ? * * 
 
 S e r v e r n   v � r d n y c k e l n   h i t t a d e s   i n t e   i   c a c h e n .   D u   h a r   i n g e n   g a r a n t i   f � r   a t t   s e r v e r n   � r   d e n   d a t o r   d u   t r o r   a t t   d e t   � r . 
 
 S e r v e r n s   % s   n y c k e l d e t a l j e r   � r : 
 
 % s 
 
 O m   d u   l i t a r   p �   d e n   h � r   v � r d e n ,   t r y c k   p �   J a .   O m   d u   v i l l   a n s l u t a   u t a n   a t t   l � g g a   t i l l   v � r d n y c k e l   i   c a c h e n   t r y c k e r   d u   p �   N e j .   F � r   a t t   a v b r y t a   a n s l u t n i n g e n   t r y c k e r   d u   p �   A v b r y t . * * V A R N I N G   -   P O T E N T I E L L T   S � K E R H E T S I N T R � N G ! * * 
 
 S e r v e r n s   v � r d n y c k e l   m a t c h a r   i n t e   d e n   s o m   W i n S C P   h a r   i   c a c h e n .   D e t   b e t y d e r   a t t   a n t i n g e n   s e r v e r n s   a d m i n i s t r a t � r   h a r   � n d r a t   v � r d n y c k e l n ,   s e r v e r n   v i s a r   o l i k a   n y c k e l a r   u n d e r   v i s s a   o m s t � n d i g h e t e r ,   e l l e r   a t t   d u   h a r   f a k t i s k t   a n s l u t i t   t i l l   e n   a n n a n   d a t o r   s o m   l � t s a s   v a r a   s e r v e r n . 
 
 N y c k l a r n a   f � r   % s   � r : 
 
 % s 
 
 O m   d u   f � r v � n t a d e   d i g   d e n n a   � n d r i n g ,   l i t a r   p �   d e n   n y a   n y c k e l n   o c h   v i l l   f o r t s � t t a   a t t   a n s l u t a   t i l l   s e r v e r n ,   t r y c k   a n t i n g e n   p �   U p p d a t e r a   f � r   a t t   u p p d a t e r a   c a c h e n   e l l e r   t r y c k   p �   L � g g   t i l l   f � r   a t t   l � g g a   t i l l   d e n   n y a   n y c k e l n   i   c a c h e n   m e d a n   d u   b e h � l l e r   d e n   g a m l a .   O m   d u   v i l l   f o r t s � t t a   a t t   a n s l u t a   m e n   u t a n   a t t   u p p d a t e r a   c a c h e n ,   t r y c k   p �   H o p p a   � v e r .   F � r   a t t   � v e r g e   a n s l u t n i n g e n   h e l t ,   t r y c k   p �   A v b r y t .   A t t   t r y c k a   p �   A v b r y t   � r   d e t   e n d a   g a r a n t e r a d e   s � k r a   v a l e t . 0D u   l a d d a r   e n   S S H - 2   p r i v a t   n y c k e l   s o m   h a r   e t t   g a m m a l t   f i l f o r m a t .   D e t   i n n e b � r   a t t   d i n   n y c k e l f i l   i n t e   � r   h e l t   s � k e r   f � r   m a n i p u l e r i n g s f � r s � k .   V i   r e k o m m e n d e r a r   d i g   a t t   k o n v e r t e r a   d i n   n y c k e l   t i l l   d e t   n y a   f o r m a t e t . 
 
 D u   k a n   u t f � r a   d e n   h � r   k o n v e r t e r i n g e n   g e n o m   a t t   l a d d a   f i l e n   i   P u T T Y g e n   o c h   s e d a n   s p a r a   d e n   i g e n . � H e l p   [   < k o m m a n d o >   [   < k o m m a n d o 2 >   . . .   ] 
     V i s a r   l i s t a   p �   k o m m a n d o n   o m   i n g a   p a r a m e t e r a r   a n g e s . 
     V i s a r   h j � l p   o m   e t t   k o m m a n d o   o m   d e t   a n g e s . 
 a l i a s : 
     m a n 
 e x e m p e l : 
     h e l p 
     h e l p   l s 
 D e x i t 
     S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t . 
 a l i a s : 
     b y e 
 o p e n   < s i t e > 
 o p e n   s f t p | s c p | f t p [ e s ] | d a v [ s ] | s 3   : / /   [   < u s e r >   [   : p a s s w o r d   ]   @   ]   < h o s t >   [   : < p o r t >   ] 
     E s t a b l i s h e s   c o n n e c t i o n   t o   g i v e n   h o s t .   U s e   e i t h e r   n a m e   o f   t h e   s i t e   o r 
     s p e c i f y   h o s t ,   u s e r n a m e ,   p o r t   a n d   p r o t o c o l   d i r e c t l y . 
 s w i t c h e s : 
     - p r i v a t e k e y = < f i l e >   S S H   p r i v a t e   k e y   f i l e 
     - h o s t k e y = < f i n g e r p r i n t >   F i n g e r p r i n t   o f   s e r v e r   h o s t   k e y   ( S F T P   a n d   S C P   o n l y ) . 
     - c l i e n t c e r t = < f i l e >   T L S / S S L   c l i e n t   c e r t i f i c a t e   f i l e 
     - c e r t i f i c a t e = < f i n g e r p r i n t >   F i n g e r p r i n t   o f   T L S / S S L   c e r t i f i c a t e 
                                           ( F T P S   a n d   W e b D A V S   o n l y ) 
     - p a s s p h r a s e = < p h r >     P r i v a t e   k e y   p a s s p h r a s e 
     - p a s s i v e = o n | o f f         P a s s i v e   m o d e   ( F T P   p r o t o c o l   o n l y ) 
     - i m p l i c i t                     I m p l i c i t   T L S / S S L   ( F T P   p r o t o c o l   o n l y ) 
     - e x p l i c i t                     E x p l i c i t   T L S / S S L   ( F T P   p r o t o c o l   o n l y ) 
     - t i m e o u t = < s e c >           S e r v e r   r e s p o n s e   t i m e o u t 
     - u s e r n a m e = < u s e r >       A n   a l t e r n a t i v e   w a y   t o   p r o v i d e   a   u s e r n a m e 
     - p a s s w o r d = < p a s s w o r d >   A n   a l t e r n a t i v e   w a y   t o   p r o v i d e   a   p a s s w o r d 
     - r a w s e t t i n g s   s e t t i n g 1 = v a l u e 1   s e t t i n g 2 = v a l u e 2   . . . 
                                           C o n f i g u r e s   a n y   s i t e   s e t t i n g s   u s i n g   r a w   f o r m a t 
                                           a s   i n   a n   I N I   f i l e 
     - f i l e z i l l a                   L o a d   < s i t e >   f r o m   F i l e Z i l l a   s i t e   m a n a g e r 
     - n e w p a s s w o r d = < p a s s w o r d >   C h a n g e s   p a s s w o r d   t o   < p a s s w o r d > 
 e x a m p l e s : 
     o p e n 
     o p e n   s f t p : / / m a r t i n @ e x a m p l e . c o m : 2 2 2 2   - p r i v a t e k e y = m y k e y . p p k 
     o p e n   m a r t i n @ e x a m p l e . c o m 
     o p e n   e x a m p l e . c o m 
 � c l o s e   [   < s e s s i o n >   ] 
     S t � n g e r   s e s s i o n   s p e c i f i c e r a d   m e d   s i t t   n u m m e r .   O m   s e s s i o n s n u m r e t   i n t e   � r 
     s p e c i f i c e r a d ,   s t � n g s   d e n   a k t u e l l a   s e s s i o n e n . 
 e x e m p e l : 
     c l o s e 
     c l o s e   1 
 � s e s s i o n   [   < s e s s i o n >   ] 
     G � r   s e s s i o n e n   s p e c i f i c e r a d   m e d   e t t   n u m m e r   a k t i v .   O m   e t t   s e s s i o n s n u m m e r 
     i n t e   � r   s p e c i f i c e r a d ,   l i s t a s   a n s l u t n a   s e s s i o n e r . 
 e x e m p e l : 
     s e s s i o n 
     s e s s i o n   1 
 ; p w d 
     V i s a r   a k t u e l l   f j � r r k a t a l o g   f � r   d e n   a k t i v a   s e s s i o n e n . 
 � c d   [   < k a t a l o g >   ] 
     � n d r a r   a k t u e l l   k a t a l o g   p �   s e r v e r n   i   d e n   a k t i v a   s e s s i o n e n . 
     O m   e n   k a t a l o g   i n t e   a n g e s ,   a n v � n d s   h e m k a t a l o g e n . 
 e x e m p e l : 
     c d   / h o m e / m a r t i n 
     c d 
 Ul s   [   < d i r e c t o r y >   ] / [   < w i l d c a r d >   ] 
     L i s t s   t h e   c o n t e n t s   o f   s p e c i f i e d   r e m o t e   d i r e c t o r y .   I f   d i r e c t o r y   i s   
     n o t   s p e c i f i e d ,   l i s t s   w o r k i n g   d i r e c t o r y . 
     W h e n   w i l d c a r d   i s   s p e c i f i e d ,   i t   i s   t r e a t e d   a s   s e t   o f   f i l e s   t o   l i s t . 
     O t h e r w i s e ,   a l l   f i l e s   a r e   l i s t e d . 
 a l i a s : 
     d i r 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     l s 
     l s   * . h t m l 
     l s   / h o m e / m a r t i n 
 @ l p w d 
     V i s a r   a k t u e l l   l o k a l   k a t a l o g   ( g � l l e r   f � r   a l l a   s e s s i o n e r ) . 
 J l c d   < k a t a l o g > 
     B y t e r   l o k a l   k a t a l o g   f � r   a l l a   s e s s i o n e r . 
 e x e m p e l : 
     c d   d : \ 
 Bl l s   [   < d i r e c t o r y >   ] \ [   < w i l d c a r d >   ] 
     L i s t s   t h e   c o n t e n t s   o f   s p e c i f i e d   l o c a l   d i r e c t o r y .   I f   d i r e c t o r y   i s   
     n o t   s p e c i f i e d ,   l i s t s   w o r k i n g   d i r e c t o r y . 
     W h e n   w i l d c a r d   i s   s p e c i f i e d ,   i t   i s   t r e a t e d   a s   s e t   o f   f i l e s   t o   l i s t . 
     O t h e r w i s e ,   a l l   f i l e s   a r e   l i s t e d . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     l l s 
     l l s   * . h t m l 
     l l s   d : \ 
 9r m   < f i l e >   [   < f i l e 2 >   . . .   ] 
     R e m o v e s   o n e   o r   m o r e   r e m o t e   f i l e s .   I f   r e m o t e   r e c y c l e   b i n   i s 
     c o n f i g u r e d ,   m o v e s   f i l e   t o   t h e   b i n   i n s t e a d   o f   d e l e t i n g   i t . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     r m   i n d e x . h t m l 
     r m   i n d e x . h t m l   a b o u t . h t m l 
     r m   * . h t m l 
 � r m d i r   < k a t a l o g >   [   < k a t a l o g 2 >   . . .   ] 
     R a d e r a r   e n   e l l e r   f l e r a   f j � r r k a t a l o g e r .   O m   f j � r r p a p p e r s k o r g e n   � r 
   k o n f i g u r e r a d ,   f l y t t a s   k a t a l o g e n   d i t   i s t � l l e t   f � r   a t t   r a d e r a s . 
 e x e m p e l : 
     r m d i r   p u b l i c _ h t m l 
 ?m v   < f i l e >   [   < f i l e 2 >   . . .   ]   [   < d i r e c t o r y > /   ] [   < n e w n a m e >   ] 
     M o v e s   o r   r e n a m e s   o n e   o r   m o r e   r e m o t e   f i l e s .   D e s t i n a t i o n   d i r e c t o r y   o r   n e w 
     n a m e   o r   b o t h   m u s t   b e   s p e c i f i e d .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h   
     s l a s h .   O p e r a t i o n   m a s k   c a n   b e   u s e d   i n s t e a d   o f   n e w   n a m e . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 a l i a s : 
     r e n a m e 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     m v   i n d e x . h t m l   p u b l i c _ h t m l / 
     m v   i n d e x . h t m l   a b o u t . * 
     m v   i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . * 
     m v   p u b l i c _ h t m l / i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . h t m l   / h o m e / m a r t i n / * . b a k 
     m v   * . h t m l   / h o m e / b a c k u p / * . b a k 
 ^c h m o d   < m o d e >   < f i l e >   [   < f i l e 2 >   . . .   ] 
     C h a n g e s   p e r m i s s i o n s   o f   o n e   o r   m o r e   r e m o t e   f i l e s .   M o d e   c a n   b e   s p e c i f i e d 
     a s   t h r e e   o r   f o u r - d i g i t   o c t a l   n u m b e r . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     c h m o d   6 4 4   i n d e x . h t m l   a b o u t . h t m l 
     c h m o d   1 7 0 0   / h o m e / m a r t i n / p u b l i c _ h t m l 
     c h m o d   6 4 4   * . h t m l 
 t l n   < m � l >   < s y m b o l i s k   l � n k > 
     S k a p a r   s y m b o l i s k   f j � r r l � n k . 
 a l i a s : 
     s y m l i n k 
 e x e m p e l : 
     l n   / h o m e / m a r t i n / p u b l i c _ h t m l   w w w 
 D m k d i r   < k a t a l o g > 
     S k a p a r   f j � r r k a t a l o g . 
 e x e m p e l : 
     m k d i r   p u b l i c _ h t m l 
 g e t   < f i l e >   [   [   < f i l e 2 >   . . .   ]   < d i r e c t o r y > \ [   < n e w n a m e >   ]   ] 
     D o w n l o a d s   o n e   o r   m o r e   f i l e s   f r o m   r e m o t e   d i r e c t o r y   t o   l o c a l   d i r e c t o r y . 
     I f   o n l y   o n e   p a r a m e t e r   i s   s p e c i f i e d   d o w n l o a d s   t h e   f i l e   t o   l o c a l   w o r k i n g 
     d i r e c t o r y .   I f   m o r e   p a r a m e t e r s   a r e   s p e c i f i e d ,   a l l   e x c e p t   t h e   l a s t   o n e 
     s p e c i f y   s e t   o f   f i l e s   t o   d o w n l o a d .   T h e   l a s t   p a r a m e t e r   s p e c i f i e s   t a r g e t 
     l o c a l   d i r e c t o r y   a n d   o p t i o n a l l y   o p e r a t i o n   m a s k   t o   s t o r e   f i l e ( s )   u n d e r 
     d i f f e r e n t   n a m e .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h   b a c k s l a s h .   
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
     T o   d o w n l o a d   m o r e   f i l e s   t o   c u r r e n t   w o r k i n g   d i r e c t o r y   u s e   ' . \ '   a s   t h e 
     l a s t   p a r a m e t e r . 
 a l i a s : 
     r e c v ,   m g e t 
 s w i t c h e s : 
     - d e l e t e                     D e l e t e   s o u r c e   r e m o t e   f i l e ( s )   a f t e r   t r a n s f e r 
     - r e s u m e                     R e s u m e   t r a n s f e r   i f   p o s s i b l e   ( S F T P   a n d   F T P   p r o t o c o l s   o n l y ) 
     - a p p e n d                     A p p e n d   f i l e   t o   e n d   o f   t a r g e t   f i l e   ( S F T P   p r o t o c o l   o n l y ) 
     - p r e s e r v e t i m e         P r e s e r v e   t i m e s t a m p 
     - n o p r e s e r v e t i m e     D o   n o t   p r e s e r v e   t i m e s t a m p 
     - s p e e d = < k b p s >         L i m i t   t r a n s f e r   s p e e d   ( i n   K B / s ) 
     - t r a n s f e r = < m o d e >   T r a n s f e r   m o d e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >   S e t s   f i l e   m a s k . 
     - r e s u m e s u p p o r t = < s t a t e >   C o n f i g u r e s   r e s u m e   s u p p o r t . 
                                       P o s s i b l e   v a l u e s   a r e   ' o n ' ,   ' o f f '   o r   t h r e s h o l d 
     - n e w e r o n l y               T r a n s f e r   n e w   a n d   u p d a t e d   f i l e s   o n l y 
     - l a t e s t                     T r a n s f e r   t h e   l a t e s t   f i l e   o n l y 
 e f f e c t i v e   o p t i o n s : 
     c o n f i r m ,   f a i l o n n o m a t c h ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     g e t   i n d e x . h t m l 
     g e t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . \ 
     g e t   i n d e x . h t m l   a b o u t . h t m l   d : \ w w w \ 
     g e t   p u b l i c _ h t m l / i n d e x . h t m l   d : \ w w w \ a b o u t . * 
     g e t   * . h t m l   * . p n g   d : \ w w w \ * . b a k 
 �p u t   < f i l e >   [   [   < f i l e 2 >   . . .   ]   < d i r e c t o r y > / [   < n e w n a m e >   ]   ] 
     U p l o a d s   o n e   o r   m o r e   f i l e s   f r o m   l o c a l   d i r e c t o r y   t o   r e m o t e   d i r e c t o r y . 
     I f   o n l y   o n e   p a r a m e t e r   i s   s p e c i f i e d   u p l o a d s   t h e   f i l e   t o   r e m o t e   w o r k i n g 
     d i r e c t o r y .   I f   m o r e   p a r a m e t e r s   a r e   s p e c i f i e d ,   a l l   e x c e p t   t h e   l a s t   o n e 
     s p e c i f y   s e t   o f   f i l e s   t o   u p l o a d .   T h e   l a s t   p a r a m e t e r   s p e c i f i e s   t a r g e t 
     r e m o t e   d i r e c t o r y   a n d   o p t i o n a l l y   o p e r a t i o n   m a s k   t o   s t o r e   f i l e ( s )   u n d e r 
     d i f f e r e n t   n a m e .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h   s l a s h .   
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
     T o   u p l o a d   m o r e   f i l e s   t o   c u r r e n t   w o r k i n g   d i r e c t o r y   u s e   ' . / '   a s   t h e 
     l a s t   p a r a m e t e r . 
 a l i a s : 
     s e n d ,   m p u t 
 s w i t c h e s : 
     - d e l e t e                           D e l e t e   s o u r c e   l o c a l   f i l e ( s )   a f t e r   t r a n s f e r 
     - r e s u m e                           R e s u m e   t r a n s f e r   i f   p o s s i b l e   ( S F T P   a n d   F T P   p r o t o c o l s   o n l y ) 
     - a p p e n d                           A p p e n d   f i l e   t o   e n d   o f   t a r g e t   f i l e   ( S F T P   p r o t o c o l   o n l y ) 
     - p r e s e r v e t i m e               P r e s e r v e   t i m e s t a m p 
     - n o p r e s e r v e t i m e           D o   n o t   p r e s e r v e   t i m e s t a m p 
     - p e r m i s s i o n s = < m o d e >   S e t   p e r m i s s i o n s 
     - n o p e r m i s s i o n s             K e e p   d e f a u l t   p e r m i s s i o n s 
     - s p e e d = < k b p s >               L i m i t   t r a n s f e r   s p e e d   ( i n   K B / s ) 
     - t r a n s f e r = < m o d e >         T r a n s f e r   m o d e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >         S e t s   f i l e   m a s k . 
     - r e s u m e s u p p o r t = < s t a t e >   C o n f i g u r e s   r e s u m e   s u p p o r t . 
                                             P o s s i b l e   v a l u e s   a r e   ' o n ' ,   ' o f f '   o r   t h r e s h o l d 
     - n e w e r o n l y                     T r a n s f e r   n e w   a n d   u p d a t e d   f i l e s   o n l y 
     - l a t e s t                           T r a n s f e r   t h e   l a t e s t   f i l e   o n l y 
 e f f e c t i v e   o p t i o n s : 
     c o n f i r m ,   f a i l o n n o m a t c h ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     p u t   i n d e x . h t m l 
     p u t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . / 
     p u t   - p e r m i s s i o n s = 6 4 4   i n d e x . h t m l   a b o u t . h t m l   / h o m e / m a r t i n / p u b l i c _ h t m l / 
     p u t   d : \ w w w \ i n d e x . h t m l   a b o u t . * 
     p u t   * . h t m l   * . p n g   / h o m e / m a r t i n / b a c k u p / * . b a k 
 �o p t i o n   [   < o p t i o n >   [   < v a l u e >   ]   ] 
     I f   n o   p a r a m e t e r s   a r e   s p e c i f i e d ,   l i s t s   a l l   s c r i p t   o p t i o n s   a n d   t h e i r 
     v a l u e s .   W h e n   o n e   p a r a m e t e r   i s   s p e c i f i e d   o n l y ,   s h o w s   v a l u e   o f   t h e   o p t i o n . 
     W h e n   t w o   p a r a m e t e r s   a r e   s p e c i f i e d   s e t s   v a l u e   o f   t h e   o p t i o n . 
     I n i t i a l   v a l u e s   o f   s o m e   o p t i o n s   a r e   t a k e n   f r o m   a p p l i c a t i o n   c o n f i g u r a t i o n , 
     h o w e v e r   m o d i f i n g   t h e   o p t i o n s   d o e s   n o t   c h a n g e   t h e   a p p l i c a t i o n 
     c o n f i g u r a t i o n . 
 o p t i o n s   a r e : 
     e c h o           o n | o f f 
                       T o g g l e s   e c h o i n g   o f   c o m m a n d   b e i n g   e x e c u t e d . 
                       C o m m a n d s   a f f e c t e d :   a l l 
     b a t c h         o n | o f f | a b o r t | c o n t i n u e 
                       T o g g l e s   b a t c h   m o d e   ( a l l   p r o m p t s   a r e   a u t o m a t i c a l l y   r e p l i e d 
                       n e g a t i v e l y ) .   W h e n   ' o n ' ,   i t   i s   r e c o m m e n d e d   t o   s e t   ' c o n f i r m ' 
                       t o   ' o f f '   t o   a l l o w   o v e r w r i t e s .   W i t h   ' a b o r t ' ,   s c r i p t   i s   a b o r t e d 
                       w h e n   a n y   e r r o r   o c c u r s .   W i t h   ' c o n t i n u e ' ,   a l l   e r r o r s   a r e   i g n o r e d . 
                       R e c o n n e c t   t i m e   i s   a u t o m a t i c a l l y   l i m i t e d   d o   1 2 0 s ,   i f   n o t   l i m i t e d   y e t . 
                       C o m m a n d s   a f f e c t e d :   n e a r l y   a l l 
     c o n f i r m     o n | o f f 
                       T o g g l e s   c o n f i r m a t i o n s   ( o v e r w r i t e ,   e t c . ) . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t 
     r e c o n n e c t t i m e   o f f   |   < s e c > 
                       T i m e   l i m i t   i n   s e c o n d s   t o   t r y   r e c o n n e c t i n g   b r o k e n   s e s s i o n s . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
     f a i l o n n o m a t c h   o n | o f f 
                       W h e n   ' o n ' ,   c o m m a n d s   f a i l   w h e n   f i l e   m a s k   m a t c h e s   n o   f i l e s . 
                       W h e n   ' o f f ' ,   c o m m a n d s   d o   n o t h i n g   w h e n   f i l e   m a s k   m a t c h e s   n o   f i l e s . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   r m ,   m v ,   c h m o d ,   l s ,   l l s 
 e x a m p l e s : 
     o p t i o n 
     o p t i o n   b a t c h 
     o p t i o n   c o n f i r m   o f f 
 As y n c h r o n i z e   l o c a l | r e m o t e | b o t h   [   < l o k a l   k a t a l o g >   [   < f j � r r k a t a l o g >   ]   ] 
     N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' l o c a l '   s y n k r o n i s e r a s   l o k a l   k a t a l o g   m e d 
     f j � r r k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' r e m o t e '   s y n k r o n i s e r a s   f j � r r k a t a l o g 
     m e d   l o k a l   k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' b o t h '   s y n k r o n i s e r a s 
     k a t a l o g e r n a   m o t   v a r a n d r a . 
     N � r   k a t a l o g e r   i n t e   s p e c i f i c e r a s ,   s y n k r o n i s e r a s   a k t u e l l 
     k a t a l o g . 
     O B S :   � v e r s k r i v n i n g s b e k r � f t e l s e r   � r   a l l t i d   a v   f � r   k o m m a n d o t . 
 v � x l a r : 
     - p r e v i e w                           F � r h a n d s g r a n s k a   � n d r i n g a r ,   s y n k r o n i s e r a r   i n t e 
     - d e l e t e                             T a   b o r t   f � r � l d r a d e   f i l e r 
     - m i r r o r                             S p e g e l l � g e   ( s y n k r o n i s e r a r   f � r � l d r a d e   f i l e r   o c k s � ) . 
                                               I g n o r e r a s   m e d   ' b o t h ' . 
     - c r i t e r i a = < k r i t e r i e r >   J � m f � r e l s e k r i t e r i e r .   M � j l i g a   v � r d e n   � r   ' n o n e ' ,   ' t i m e ' , 
                                               ' s i z e '   o c h   ' e i t h e r ' .   I g n o r e r a s   m e d   ' b o t h ' - l � g e . 
     - p e r m i s s i o n s = < l � g e >     A n g e   r � t t i g h e t e r 
     - n o p e r m i s s i o n s               B e h � l l   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k b p s >               B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
     - t r a n s f e r = < l � g e >           � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >           A n g e   f i l m a s k . 
     - r e s u m e s u p p o r t = < t i l l s t � n d >   K o n f i g u r e r a r   � t e r u p p t a g n i n g s s t � d . 
                                               M � j l i g a   v � r d e n   � r   ' o n ' ,   ' o f f '   e l l e r   t r � s k e l 
 e f f e k t i v a   a l t e r n a t i v : 
     r e c o n n e c t t i m e 
 e x e m p e l : 
     s y n c h r o n i z e   r e m o t e   - d e l e t e 
     s y n c h r o n i z e   b o t h   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 Sk e e p u p t o d a t e   [   < l o c a l   d i r e c t o r y >   [   < r e m o t e   d i r e c t o r y >   ]   ] 
     W a t c h e s   f o r   c h a n g e s   i n   l o c a l   d i r e c t o r y   a n d   r e f l e c t s   t h e m   o n   r e m o t e   o n e . 
     W h e n   d i r e c t o r i e s   a r e   n o t   s p e c i f i e d ,   c u r r e n t   w o r k i n g   d i r e c t o r i e s   a r e 
     s y n c h r o n i z e d .   T o   s t o p   w a t c h i n g   f o r   c h a n g e s   p r e s s   C t r l - C . 
     N o t e :   O v e r w r i t e   c o n f i r m a t i o n s   a r e   a l w a y s   o f f   f o r   t h e   c o m m a n d . 
 s w i t c h e s : 
     - d e l e t e                           D e l e t e   o b s o l e t e   f i l e s 
     - p e r m i s s i o n s = < m o d e >   S e t   p e r m i s s i o n s 
     - n o p e r m i s s i o n s             K e e p   d e f a u l t   p e r m i s s i o n s 
     - s p e e d = < k b p s >               L i m i t   t r a n s f e r   s p e e d   ( i n   K B / s ) 
     - t r a n s f e r = < m o d e >         T r a n s f e r   m o d e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >         S e t s   f i l e   m a s k . 
     - r e s u m e s u p p o r t = < s t a t e >   C o n f i g u r e s   r e s u m e   s u p p o r t . 
                                             P o s s i b l e   v a l u e s   a r e   ' o n ' ,   ' o f f '   o r   t h r e s h o l d 
 e f f e c t i v e   o p t i o n s : 
     r e c o n n e c t t i m e 
 e x a m p l e s : 
     k e e p u p t o d a t e   - d e l e t e 
     k e e p u p t o d a t e   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 Wc a l l   < K o m m a n d o > 
     M e d   S F T P   o c h   S C P   p r o t o k o l l e n ,   k � r s   g o d t y c k l i g t   f j � r r s k a l s k o m m a n d o . 
     O m   a k t u e l l   s e s s i o n   i n t e   t i l l � t e r   k � r n i n g   a v   g o d t y c k l i g   f j � r r k o m m a n d o 
     s k i l d a   s k a l s e s s i o n e r   k o m m e r   a t t   � p p n a s   a u t o m a t i s k t . 
     O m   F T P   p r o t o k o l l ,   k � r   e t t   p r o t o k o l l k o m m a n d o . 
     K o m m a n d o t   k a n   i n t e   k r � v a   a n v � n d a r i n p u t . 
 a l i a s : 
     ! 
 e x e m p e l : 
     c a l l   t o u c h   i n d e x . h t m l 
 ] e c h o   < m e d d e l a n d e > 
     S k r i v e r   m e d d e l a n d e   t i l l   s k r i p t u t d a t a . 
 e x e m p e l : 
     e c h o   S t a r t i n g   u p l o a d . . . 
 Y s t a t   < f i l > 
     H � m t a r   o c h   l i s t a r   a t t r i b u t   f � r   a n g i v e n   f j � r r f i l . 
 e x e m p e l : 
     s t a t   i n d e x . h t m l 
 a c h e c k s u m   < a l g >   < f i l e > 
     C a l c u l a t e s   c h e c k s u m   o f   r e m o t e   f i l e . 
 e x a m p l e : 
     c h e c k s u m   s h a - 1   i n d e x . h t m l 
 (c p   < f i l e >   [   < f i l e 2 >   . . .   ]   [   < d i r e c t o r y > /   ] [   < n e w n a m e >   ] 
     D u p l i c a t e s   o n e   o r   m o r e   r e m o t e   f i l e s .   D e s t i n a t i o n   d i r e c t o r y   o r   n e w 
     n a m e   o r   b o t h   m u s t   b e   s p e c i f i e d .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h 
     s l a s h .   O p e r a t i o n   m a s k   c a n   b e   u s e d   i n s t e a d   o f   n e w   n a m e . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     c p   i n d e x . h t m l   p u b l i c _ h t m l / 
     c p   i n d e x . h t m l   a b o u t . * 
     c p   i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . * 
     c p   p u b l i c _ h t m l / i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . h t m l   / h o m e / m a r t i n / * . b a k 
     c p   * . h t m l   / h o m e / b a c k u p / * . b a k 
             
 C O R E _ E R R O R " V � r d n y c k e l n   k u n d e   i n t e   v e r i f i e r a s !  A n s l u t n i n g   m i s s l y c k a d e s .  A v s l u t a d   a v   a n v � n d a r e n .  T a p p a d   a n s l u t n i n g . # K a n   i n t e   h i t t a   k o m m a n d o t s   r e t u r k o d . C K o m m a n d o t   ' % s ' 
 m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d   o c h   f e l m e d d e l a n d e 
 % s . ) K o m m a n d o t   m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d . 7 K o m m a n d o t   ' % s '   m i s s l y c k a d e s   m e d   o g i l t i g   u t m a t n i n g   ' % s ' . = F e l   u p p s t o d   n � r   n a m n e t   p �   a k t u e l l   f j � r r k a t a l o g   s k u l l e   h � m t a s . | F e l   u p p s t o d   n � r   s t a r t m e d d e l a n d e   h o p p a d e s   � v e r .   D i t t   s k a l   � r   a n t a g l i g e n   i n k o m p a t i b e l t   m e d   a p p l i k a t i o n e n   ( B A S H   r e k o m m e n d e r a s ) . ) F e l   u p p s t o d   n � r   k a t a l o g   b y t t e s   t i l l   ' % s ' .     ) F e l   u p p s t o d   n � r   l i s t n i n g   a v   k a t a l o g   ' % s ' . % O v � n t a d   k a t a l o g l i s t n i n g   v i d   r a d   ' % s ' . # F e l a k t i g   r � t t i g h e t s b e s k r i v n i n g   ' % s ' ; F e l   u p p s t o d   n � r   d e n   a l l m � n n a   k o n f i g u r a t i o n e n   s k u l l e   r e n s a s .   F e l   v i d   r e n s n i n g   a v   c a c h e m i n n e t . 1 F e l   u p p s t o d   n � r   f i l e n   m e d   s l u m p t a l s f r � n   r e n s a d e s . - F e l   u p p s t o d   n � r   c a c h a d e   v � r d n y c k l a r   r e n s a d e s . Q F e l   u p p s t o d   n � r   v a r i a b e l   i n n e h � l l a n d e   r e t u r k o d   a v   s e n a s t e   k o m m a n d o   s k u l l e   h i t t a s . 0 F e l   u p p s t o d   n � r   a n v � n d a r g r u p p e r   s k u l l e   s l � s   u p p . " F i l   e l l e r   k a t a l o g   ' % s '   f i n n s   i n t e . ) K a n   i n t e   h i t t a   a t t r i b u t e n   f � r   f i l e n   ' % s ' .  K a n   i n t e   � p p n a   f i l e n   ' % s ' . ( F e l   u p p s t o d   n � r   f i l e n   ' % s '   s k u l l e   l � s a s . 3 A l l v a r l i g t   f e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l e n   ' % s ' . 0 F i l k o p i e r i n g e n   t i l l   f j � r r k a t a l o g e n   m i s s l y c k a d e s .   0 F i l k o p i e r i n g e n   f r � n   f j � r r k a t a l o g e n   m i s s l y c k a d e s . % S C P   p r o t o k o l l f e l :   O v � n t a d   r a d b r y t n i n g & S C P   p r o t o k o l l f e l :   F e l a k t i g t   t i d s f o r m a t 2 S C P   p r o t o k o l l f e l :   F e l a k t i g   c o n t r o l   r e c o r d   ( % s ;   % s ) # K o p i e r i n g   a v   f i l   ' % s '   m i s s l y c k a d e s . 1 S C P   p r o t o k o l l f e l :   F e l a k t i g t   f i l b e s k r i v n i n g s f o r m a t  ' % s '   � r   i n g e n   k a t a l o g ! ( F e l   u p p s t o d   n � r   k a t a l o g e n   ' % s '   s k a p a d e s .  K a n   i n t e   s k a p a   f i l e n   ' % s ' . * F e l   u p p s t o d   v i d   s k r i v n i n g   t i l l   f i l e n   ' % s ' . * K a n   i n t e   s � t t a   a t t r i b u t e n   t i l l   f i l e n   ' % s ' . + F e l m e d d e l a n d e   m o t t a g e t   f r � n   f j � r r s i d a :   ' % s ' " F e l   v i d   b o r t t a g n i n g   a v   f i l e n   ' % s ' . 7 F e l   u p p s t o d   v i d   l o g g n i n g   o c h   d e n   h a r   d � r f � r   s t � n g t s   a v .  K a n   i n t e   � p p n a   l o g g f i l e n   ' % s ' . 0 F e l   u p p s t o d   n � r   f i l e n   ' % s '   b y t t e   n a m n   t i l l   ' % s ' .     F i l e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . $ K a t a l o g e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . 2 F e l   u p p s t o d   v i d   b y t e   a v   k a t a l o g   t i l l   h e m k a t a l o g e n . ' F e l   u p p s t o d   v i d   r e n s n i n g   a v   a l l a   a l i a s .   ; F e l   u p p s t o d   n � r   n a t i o n e l l a   a n v � n d a r v a r i a b l e r   s k u l l e   r e n s a s . ! O v � n t a d   i n d a t a   f r � n   s e r v e r n :   ' % s ' ( F e l   u p p s t o d   n � r   I N I - f i l e n   s k u l l e   r e n s a s .   6 A u t e n t i s e r i n g s l o g g   ( s e   s e s s i o n s l o g g   f � r   d e t a l j e r ) : 
 % s 
  A u t e n t i s e r i n g   m i s s l y c k a d e s . # A n s l u t n i n g e n   h a r   o v � n t a t   a v s l u t a t s . 1 F e l   u p p s t o d   n � r   n y c k e l n   s p a r a d e s   t i l l   f i l e n   ' % s ' .   ) S e r v e r n   s k i c k a d e   k o m m a n d o t   s l u t s t a t u s   % d . < S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g   m e d d e l a n d e t y p   v i d   s v a r   ( % d ) .   I S F T P - s e r v e r n s   v e r s i o n   ( % d )   s t � d s   i n t e .   V e r s i o n e r   s o m   s t � d s   � r   % d   t i l l   % d . E S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g t   m e d d e l a n d e n u m m e r   % d   ( f � r v � n t a d e   % d ) .  O v � n t a d   O K   r e s p o n s .  O v � n t a d   E O F   r e s p o n s . ! F i l e n   e l l e r   k a t a l o g e n   f i n n s   i n t e .  � t k o m s t   n e k a d . . A l l m � n t   f e l   ( s e r v e r n   b o r d e   g e   f e l b e s k r i v n i n g ) . J D � l i g t   m e d d e l a n d e   ( D � l i g t   f o r m a t e r a t   p a k e t   e l l e r   i n k o m p a t i b e l t   p r o t o k o l l ) .  I n g e n   a n s l u t n i n g .  F � r l o r a d   a n s l u t n i n g .   S e r v e r n   s t � d e r   i n t e   o p e r a t i o n e n . - % s 
 F e l k o d :   % d 
 F e l m e d d e l a n d e   f r � n   s e r v e r % s :   % s  O k � n d   s t a t u s k o d . ' F e l   v i d   l � s n i n g   a v   s y m b o l i s k   l � n k   ' % s ' . 4 S e r v e r n   r e t u r n e r a d e   t o m   l i s t n i n g   f � r   k a t a l o g e n   ' % s ' . 6 M o t t o g   S S H _ F X P _ N A M E   p a k e t   m e d   n o l l   e l l e r   f l e r a   p o s t e r .   + K a n   i n t e   f �   d e n   v e r k l i g a   s � k v � g e n   f � r   ' % s ' . ) K a n   i n t e   � n d r a   e g e n s k a p e r   f � r   f i l e n   ' % s ' . F K a n   i n t e   i n i t i a l i s e r a   S F T P - p r o t o k o l l e t .   K � r   v � r d d a t o r n   e n   S F T P - s e r v e r ? " K a n   i n t e   l � s a   t i d s z o n s i n f o r m a t i o n .  K a n   i n t e   s k a p a   f j � r r f i l   ' % s ' .  K a n   i n t e   � p p n a   f j � r r f i l   ' % s ' .  K a n   i n t e   s t � n g a   f j � r r f i l   ' % s ' .  ' % s '   � r   i n t e   e n   f i l ! � � v e r f � r i n g e n   l y c k a d e s   s l u t f � r a ,   m e n   t e m p o r � r   � v e r f � r i n g s f i l   ' % s '   k u n d e   i n t e   b y t a   n a m n   t i l l   m � l f i l   ' % s ' .   O m   p r o b l e m e t   k v a r s t � r ,   p r o v a   m e d   a t t   s l �   a v   f i l � v e r f � r i n g e n s   � t e r u p p t a - f u n k t i o n  K a n   i n t e   s k a p a   l � n k   ' % s ' .  O g i l t i g t   k o m m a n d o   ' % s ' .  I n g e n 4 ' % s '   � r   i n g e n   t i l l � t e n   f i l r � t t i g h e t   i   o k t a l t   f o r m a t . 5 S e r v e r n   k r � v e r   e t t   e j   s t � t t   s l u t - p � - r a d   s e k v e n s   ( % s ) .  O k � n d   f i l t y p   ( % d )  O g i l t i g t   v e r k t y g .   % S � k v � g e n   f i n n s   i n t e   e l l e r   � r   o g i l t i g .  F i l e n   f i n n s   r e d a n . R F i l e n   l i g g e r   p �   e n   e n h e t   s o m   e n d a s t   s t � d e r   l � s n i n g ,   e l l e r   e n h e t e n   � r   s k r i v s k y d d a d .   D e t   f i n n s   i n g e t   m e d i a   i   e n h e t e n . * F e l   u p p s t o d   v i d   a v k o d n i n g   a v   U T F - 8   s t r � n g . < F e l   u p p s t o d   v i d   k � r n i n g   a v   e g e t   k o m m a n d o   ' % s '   p �   f i l e n   ' % s ' .  K a n   i n t e   l a d d a   l o c a l e   % d . + M o t t o g   e j   k o m p l e t t a   d a t a p a k e t   f � r e   f i l s l u t . 8 F e l   u p p s t o d   v i d   b e r � k n i n g   a v   s t o r l e k   f � r   k a t a l o g e n   ' % s ' . L M o t t o g   e t t   f � r   s t o r t   ( % d   B )   S F T P   p a k e t .   M a x i m a l t   s t � d d   p a k e t s t o r l e k   � r   % d   B . � K a n   i n t e   k � r a   S C P   f � r   a t t   s t a r t a   � v e r f � r i n g .   K o n t r o l l e r a   a t t   S C P   � r   i n s t a l l e r a t   p �   s e r v e r n   o c h   a t t   s � k v � g e n   � r   i n k l u d e r a d   i   P A T H .   D u   k a n   o c k s �   p r o v a   S F T P   i s t � l l e t   f � r   S C P .  P l a t s p r o f i l e n   ' % s '   f i n n s   r e d a n . , F e l   u p p s t o d   v i d   f l y t t   a v   f i l   ' % s '   t i l l   ' % s ' . x % s 
   
 F e l e t   o r s a k a s   n o r m a l t   a v   e t t   m e d d e l a n d e   f r � n   e t t   i n l o g g n i n g s s k r i p t   ( s o m   . p r o f i l e ) .   M e d d e l a n d e t   k a n   s t a r t a   m e d   " % s " . � * * � v e r f � r i n g   a v   f i l   ' % s '   l y c k a d e s ,   m e n   f e l   u p p s t o d   v i d   i n s t � l l n i n g   a v   r � t t i g h e t e r   o c h / e l l e r   t i d s s t � m p e l . * * 
 
 O m   p r o b l e m e t   k v a r s t � r ,   s t � n g   a v   a n g e   r � t t i g h e t e r   e l l e r   b e v a r a   t i d s s t � m p e l .   A l t e r n a t i v e t   k a n   d u   a k t i v e r a   a l t e r n a t i v e t   ' I g n o r e r a   r � t t i g h e t s f e l ' .  O g i l t i g   � t k o m s t   t i l l   m i n n e t .   2 D e t   f i n n s   i n g e n   l e d i g t   u t r y m m e   k v a r   i   f i l s y s t e m e t . t O p e r a t i o n e n   k a n   i n t e   s l u t f � r a s   p �   g r u n d   a v   a t t   d e t   s k u l l e   m e d f � r a   a t t   a n v � n d a r e n s   l a g r i n g s - q u o t a   s k u l l e   � v e r s k r i d a s . $ P r i n c i p a l   ( % s )   � r   o k � n t   f � r   s e r v e r n . 0 F e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l   ' % s '   t i l l   ' % s ' . ( O a v s l u t a t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . $ O k � n t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . V K a n   i n t e   k o m b i n e r a   f i l n a m n s m � n s t e r   ( b � r j a r   v i d   % d )   m e d   f i l l i s t m � n s t e r   ( b � r j a r   v i d   % d ) .  O k � n t   k o m m a n d o   ' % s ' . 0 T v e t y d i g t   k o m m a n d o   ' % s ' .   M � j l i g   m a t c h n i n g   � r :   % s $ P a r a m e t e r   s a k n a s   f � r   k o m m a n d o t   ' % s ' . ( F � r   m � n g a   p a r a m e t r a r   f � r   k o m m a n d o t   ' % s ' .          I n g e n   s e s s i o n .  O g i l t i g t   s e s s i o n s n u m m e r   ' % s ' .  O k � n t   a l t e r n a t i v   ' % s ' . % O k � n t   v � r d e   ' % s '   f � r   a l t e r n a t i v   ' % s ' . ( K a n   i n t e   b e s t � m m a   s t a t u s   p �   s o c k e t   ( % d ) . � F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' .   E f t e r   � t e r u p p t a g e n   f i l � v e r f � r i n g   m � s t e   b e f i n t l i g   m � l f i l   t a s   b o r t .   O m   d u   i n t e   h a   r � t t i g h e t e r   a t t   t a   b o r t   m � l f i l ,   m � s t e   d u   a v a k t i v e r a   � t e r u p p t a g n i n g   a v   f i l � v e r f � r i n g . 5 F e l   u p p s t o d   v i d   a v k o d n i n g   a v   S F T P   p a k e t   ( % d ,   % d ,   % d ) . 1 O g i l t i g t   n a m n   ' % s ' .   N a m n   k a n   i n t e   i n n e h � l l a   ' % s ' . @ F i l e n   k u n d e   i n t e   � p p n a s   f � r   a t t   d e n   � r   l � s t   a v   e n   a n n a n   p r o c e s s .  K a t a l o g e n   � r   i n t e   t o m . + D e n   s p e c i f i c e r a d e   f i l e n   � r   i n t e   e n   k a t a l o g .  F i l n a m n e t   � r   i n t e   g i l t i g t . ( F � r   m � n g a   s y m b o l i s k a   l � n k a r   a n t r � f f a d e s .  F i l e n   k a n   i n t e   t a s   b o r t . p E n   a v   p a r a m e t r a r n a   v a r   u t a n f � r   i n t e r v a l l e t ,   e l l e r   p a r a m e t r a r n a   s o m   s p e c i f i c e r a d e s   k a n   i n t e   a n v � n d a s   t i l l s a m m a n s . V D e n   s p e c i f i c e r a d e   f i l e n   v a r   e n   k a t a l o g ,   i   e n   k o n t e x t   d � r   e n   k a t a l o g   i n t e   k a n   a n v � n d a s .  L � s   f � r   b y t e i n t e r v a l l   k r o c k a d e .    L � s   f � r   b y t e i n t e r v a l l   n e k a d e s . P E n   o p e r a t i o n   f � r s � k t e   g � r a s   p �   e n   f i l   s o m   h a r   e n   v � n t a n d e   b o r t t a g n i n g s o p e r a t i o n . F F i l e n   � r   k o r r u p t ;   e n   k o n t r o l l   a v   i n t e g r i t e t e n   i   f i l s y s t e m e t   b � r   k � r a s . ? F i l   ' % s '   i n n e h � l l e r   i n t e   d e n   p r i v a t a   n y c k e l n   i   e t t   k � n t   f o r m a t . e * * D e n   p r i v a t a   n y c k e l f i l e n   ' % s '   i n n e h � l l e r   n y c k e l n   i   f o r m a t e t   % s .   W i n S C P   s t � d e r   e n d a s t   P u T T Y - f o r m a t . * * i P r i v a t   n y c k e l f i l   ' % s '   i n n e h � l l e r   n y c k e l   i   % s   f o r m a t .   D e n   f � l j e r   i n t e   d i n   f � r e d r a g n a   S S H   p r o t o k o l l v e r s i o n . � K a n   i n t e   s k r i v a   � v e r   f j � r r f i l e n   ' % s ' . $ $ 
 
 T r y c k   ' T a   b o r t '   f � r   a t t   t a   b o r t   f i l e n   o c h   s k a p a   e n   n y   i   s t � l l e t   f � r   a t t   s k r i v a   � v e r   d e n . $ $  & T a   b o r t = F e l   u p p s t o d   v i d   k o n t r o l l   a v   l e d i g t   u t r y m m e   f � r   s � k v � g e n   ' % s ' . S K a n   i n t e   h i t t a   l e d i g   l o k a l   l i s t n i n g s p o r t n u m m e r   f � r   t u n n e l   i   i n t e r v a l l e t   % d   t i l l   % d . * K a n   i n t e   u t f � r a   n � t v e r k s h � n d e l s e   ( f e l   % d ) . / S e r v e r n   a v s l u t a d e   o v � n t a t   n � t v e r k s a n s l u t n i n g e n . 1 F e l   u p p s t o d   n � r   a n s l u t n i n g e n   s k u l l e   t u n n l a s . 
   
 % s 9 F e l   u p p s t o d   n � r   k o n t r o l l s u m m a n   b e r � k n a d e s   f � r   f i l e n   ' % s ' .  I n t e r n t   f e l   % s   ( % s ) .  O p e r a t i o n e n   s t � d s   i n t e .  � t k o m s t   n e k a d . ' F r � g a r   e f t e r   a u t e n t i s e r i n g s u p p g i f t e r . . . $ O g i l t i g t   s v a r   t i l l   % s   k o m m a n d o   ' % s ' .    O k � n d   v � x e l   ' % s ' . ) F e l   u p p s t o d   v i d   � v e r f � r i n g   a v   f i l e n   ' % s ' .  K a n   i n t e   k � r a   ' % s ' .  F i l e n   ' % s '   h i t t a d e s   i n t e . . E t t   f e l   u p p s t o d   n � r   d o k u m e n t e t   s k u l l e   s t � n g a s . % ' % s '   � r   i n g e n   g i l t i g   h a s t i g h e t s g r � n s .  C e r t i f i k a t k e d j a n   � r   f � r   l � n g .  C e r t i f i k a t   h a r   u p p h � r t .   C e r t i f i k a t   � r   � n n u   i n t e   g i l t i g t .  C e r t i f i k a t   a v v i s a t .  C e r t i f i k a t   s i g n a t u r f e l .  C e r t i f i k a t   e j   s � k e r t .    S j � l v s i g n e r a t   c e r t i f i k a t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - t i l l   f � l t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - f r � n   f � l t .  O g i l t i g   C A   c e r t i f i k a t .  E j   s t � t t   c e r t i f i k a t   � n d a m � l . 5 N y c k e l a n v � n d n i n g   i n k l u d e r a r   i n t e   c e r t i f i k a t s i g n e r i n g . , B e g r � n s n i n g a r   f � r   s � k v � g s l � n g d e n   � v e r s k r i d s . + S j � l v s i g n e r a t   c e r t i f i k a t   i   c e r t i f i k a t k e d j a . 6 D e t   g � r   i n t e   a t t   a v k o d a   u t f � r d a r e n s   o f f e n t l i g a   n y c k e l . 3 D e t   g � r   i n t e   a t t   d e k r y p t e r a   c e r t i f i k a t e t s   s i g n a t u r . + D e t   g � r   i n t e   a t t   f �   u t f � r d a r e n s   c e r t i f i k a t . 2 D e t   g � r   i n t e   a t t   h � m t a   l o k a l t   u t f � r d a t   c e r t i f i k a t . 3 D e t   g � r   i n t e   a t t   v e r i f i e r a   d e t   f � r s t a   c e r t i f i k a t e t . % O k � n t   f e l   v i d   k o n t r o l l   a v   c e r t i f i k a t . 6 F e l e t   i n t r � f f a d e   p �   e t t   d j u p   a v   % d   i   c e r t i f i k a t k e d j a n .      M a s k e n   � r   o g i l t i g   n � r a   ' % s ' . � S e r v e r n   k a n   i n t e   � p p n a   a n s l u t n i n g   i   a k t i v t   l � g e .   O m   d u   s i t t e r   b a k o m   e n   N A T - r o u t e r ,   k a n   d u   b e h � v a   a n g e   e n   e x t e r n   I P - a d r e s s .   A l t e r n a t i v t ,   � v e r v � g a   a t t   b y t a   t i l l   p a s s i v t   l � g e . ( F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' . ? O g i l t i g t   v � r d e   p �   v � x e l   ' % s ' .   G i l t i g a   v � r d e n   � r   ' o n '   o c h   ' o f f ' .   0 K a n   i n t e   � p p n a   w e b b p l a t s k a t a l o g   e l l e r   a r b e t s y t a . ) N � t v e r k s f e l :   I n g e   v � g   t i l l   v � r d   " % H O S T % " . 2 N � t v e r k s f e l :   M j u k v a r a   o r s a k a d e   a v b r u t e n   a n s l u t n i n g  V � r d   " % H O S T % "   f i n n s   i n t e . 0 I n k o m m a n d e   p a k e t   v a r   f � r v a n s k a t   v i d   d e k r y p t e r i n g U % s 
 
 H j � l p   o s s   a t t   f � r b � t t r a   W i n S C P   g e n o m   a t t   r a p p o r t e r a   f e l   p �   W i n S C P : s   s u p p o r t f o r u m . - F e l   v i d   a v k o d n i n g   a v   T L S / S S L - c e r t i f i k a t   ( % s ) .  C O R E _ C O N F I R M A T I O N M V � r d e n   k o m m u n i c e r a r   i n t e   u n d e r   % d   s e k u n d e r . 
 
 V � n t a   y t t e r l i g a r e   % 0 : d   s e k u n d e r ?    & L � s e n o r d   f � r   n y c k e l n   ' % s ' : # F i l e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ' K a t a l o g e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? � D e n   f � r s t a   % s   s o m   s t � d s   a v   s e r v e r n   � r   % s ,   s o m   l i g g e r   u n d e r   d e t   k o n f i g u r e r a d e   v a r n i n g s g r � n s e n . 
 
 V i l l   d u   f o r t s � t t a   m e d   d e n   h � r   a n s l u t n i n g e n ?  c h i f f e r  k l i e n t - t i l l - s e r v e r   c h i f f e r  s e r v e r - t i l l - k l i e n t   c h i f f e r � * * V i l l   d u   � t e r u p p t a   f i l � v e r f � r i n g e n ? * * 
 
 M � l k a t a l o g e n   i n n e h � l l e r   d e l v i s   � v e r f � r d   f i l   ' % s ' . 
 
 O B S : S v a r a   ' N e j '   t a r   b o r t   d e l v i s   � v e r f � r d   f i l   o c h   s t a r t a r   o m   � v e r f � r i n g . o M � l k a t a l o g e n   i n n e h � l l e r   d e n   d e l v i s   � v e r f � r d a   f i l e n   ' % s ' ,   s o m   � r   s t � r r e   � n   k � l l f i l e n .   F i l e n   k o m m e r   a t t   t a s   b o r t . u * * V i l l   d u   l � g g a   t i l l   f i l e n   ' % s '   i   s l u t e t   a v   b e f i n t l i g   f i l ? * * 
 
 T r y c k   ' N e j '   f � r   a t t   � t e r u p p t a   f i l � v e r f � r i n g e n   i s t � l l e t . 4 % s 
   
 N y :             	 % s   b y t e s ,   % s 
 B e f i n t l i g :   	 % s   b y t e s ,   % s ' F i l e n   ' % s '   � r   s k r i v s k y d d a d .   S k r i v   � v e r ? � * * S k r i v   � v e r   l o k a l   f i l   ' % s ' ? * * M � l k a t a l o g e n   i n n e h � l l e r   r e d a n   f i l e n   ' % s ' . 
 V � l j   o m   d u   v i l l   s k r i v a   � v e r   f i l e n   e l l e r   h o p p a   � v e r   d e n n a   � v e r f � r i n g   o c h   b e h � l l a   b e f i n t l i g   f i l . � * * S k r i v   � v e r   f j � r r f i l   ' % s ' ? * * M � l k a t a l o g e n   i n n e h � l l e r   r e d a n   f i l e n   ' % s ' . 
 V � l j   o m   d u   v i l l   s k r i v a   � v e r   f i l e n   e l l e r   h o p p a   � v e r   d e n n a   � v e r f � r i n g   o c h   b e h � l l a   b e f i n t l i g   f i l .           � V � r d   k o m m u n i c e r a r   i n t e   m e r   � n   n � g r a   ' % d '   s e k u n d e r .   V � n t a r   f o r t f a r a n d e . . . 
 
 O B S :   O m   p r o b l e m e t   u p p r e p a s ,   p r o v a   a t t   s t � n g a   a v   ' O p t i m e r a   s t o r l e k e n   p �   a n s l u t n i n g s b u f f e r t ' .    & � t e r a n s l u t 
 N y t t   n a & m n      T u n n e l   f � r   % s  L � s e n o r d  L � s e n o r d   f � r   n y c k e l  S e r v e r p r o m p t  A n v � n d a r n a m n  A & n v � n d a r n a m n :  S e r v e r p r o m p t :   % s  N y t t   l � s e n o r d  S & v a r :    A n v � n d e r   T I S   a u t e n t i s e r i n g . % s $ A n v � n d e r   K r y p t o k o r t   a u t e n t i s e r i n g . % s 
 & L � s e n o r d : 0 A n v � n d e r   t a n g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % s  N & u v a r a n d e   l � s e n o r d :  & N y t t   l � s e n o r d  & B e k r � f t a   n y t t   l � s e n o r d :  A u t e n t i s e r a r   t u n n e l   g e n o m   % s  � v e r f � r   m e d   e t t   a n n a t   n a m n  & N y t t   n a m n : g* * S e r v e r n s   c e r t i f i k a t   � r   i n t e   k � n t .   D u   h a r   i n g e n   g a r a n t i   f � r   a t t   s e r v e r n   � r   d e n   d a t o r   s o m   d u   t r o r   a t t   d e   � r . * * 
 
 S e r v e r c e r t i f i k a t e t s   d e t a l j e r   f � l j e r : 
 
 % s 
 
 O m   d u   l i t a r   p �   c e r t i f i k a t e t ,   t r y c k   p �   ' J a ' .   F � r   a t t   a n s l u t a   u t a n   a t t   l a g r a   c e r t i f i k a t   t r y c k e r   d u   p �   ' N e j ' .   F � r   a t t   a v b r y t a   a n s l u t n i n g e n   t r y c k e r   p �   A v b r y t . 
 
 V i l l   d u   f o r t s � t t a   a n s l u t a   o c h   l a g r a   c e r t i f i k a t e t ? - -   O r g a n i s a t i o n :   % s 
 | -   P l a t s :   % s 
 | -   A n n a t :   % s 
  % s ,   % s c U t g i v a r e : 
 % s 
 � m n e : 
 % s 
 G i l t i g :   % s   -   % s 
 
 F i n g e r a v t r y c k : 
 -   S H A - 2 5 6 :   % s 
 -   S H A - 1 :   % s 
 
 S a m m a n f a t t n i n g :   % s $ & L � s e n o r d s f r a s   f � r   k l i e n t c e r t i f i k a t : " L � s e n o r d s f r a s   f � r   k l i e n t c e r t i f i k a t   E * * V i l l   d u   k o n v e r t e r a   d e n n a   % s   p r i v a t a   n y c k e l   t i l l   P u T T Y   f o r m a t ? * * 
 
 % s * * � r   d u   s � k e r   p �   a t t   d u   v i l l   � v e r f � r a   f l e r a   f i l e r   t i l l   e n   e n d a   f i l   ' % s '   i   e n   k a t a l o g   ' % s ' ? * * 
 
 F i l e r   k o m m e r   a t t   s k r i v a s   � v e r . 
 
 O m   d u   v e r k l i g e n   v i l l   � v e r f � r a   a l l a   f i l e r   t i l l   e n   k a t a l o g   ' % s ' ,   b e h � l l a   d e r a s   n a m n ,   s e   t i l l   a t t   d u   a v s l u t a r   s � k v � g e n   m e d   e t t   s n e d s t r e c k .  n y c k e l b y t e s a l g o r i t m  v � r d n y c k e l t y p  � t k o m s t n y c k e l - I D  � & t k o m s t n y c k e l - I D :  H e m l i g   � t k o m s t n y c k e l  H e m l i g   � t k o m s t & n y c k e l : [ D i r e k t   d u b b l e r i n g   a v   m a p p a r   s t � d s   i n t e .   A n v � n d   e n   d u b b l e r i n g   v i a   e n   l o k a l   t i l l f � l l i g   k o p i a .  A n g e   m � l   f � r   t e m p o r � r   l a g r i n g .                C O R E _ I N F O R M A T I O N  J a  N e j G V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 P r i v a t   n y c k e l f i l :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s  V e r s i o n   % s   ( % s ) > O p e r a t i o n e n   s l u t f � r d e s   f r a m g � n g s r i k t .   A n s l u t n i n g e n   a v s l u t a d e s .  S F T P - % d : S F T P   p r o t o k o l l e t s   v e r s i o n   t i l l � t e r   i n t e   n a m n b y t e   p �   f i l e r . ' S e r v e r n   s t � d e r   i n g a   u t � k n i n g a r   a v   S F T P . ( S e r v e r n   s t � d e r   f � l j a n d e   S F T P   u t � k n i n g a r :     
 L � & g g   t i l l  E n d a s t   n & y a r e  V i s a r   h j � l p . S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t    A n s l u t e r   t i l l   s e r v e r  S t � n g e r   s e s s i o n e n 4 L i s t a r   a n s l u t n a   s e s s i o n e r   e l l e r   v � l j e r   a k t i v   s e s s i o n  V i s a r   a k t u e l l   f j � r r k a t a l o g  B y t e r   a k t u e l l   f j � r r k a t a l o g  V i s a r   i n n e h � l l e t   i   f j � r r k a t a l o g  V i s a r   a k t u e l l   l o k a l   k a t a l o g  B y t e r   a k t u e l l   l o k a l   k a t a l o g ! L i s t a r   i n n e h � l l e t   i   l o k a l   k a t a l o g  T a r   b o r t   f j � r r f i l  T a r   b o r t   f j � r r k a t a l o g $ F l y t t a r   e l l e r   b y t e r   n a m n   p �   f j � r r f i l   � n d r a r   r � t t i g h e t e r n a   p �   f j � r r f i l  S k a p a r   e n   s y m b o l i s k   f j � r r l � n k  S k a p a r   f j � r r k a t a l o g 3 L a d d a r   n e r   f i l   f r � n   f j � r r k a t a l o g   t i l l   l o k a l   k a t a l o g 3 L a d d a r   u p p   f i l   f r � n   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g - S � t t e r   e l l e r   v i s a r   v � r d e n   p �   s c r i p t a l t e r n a t i v , S y n k r o n i s e r a r   f j � r r k a t a l o g   m e d   l o k a l   k a t a l o g D K o n t i n u e r l i g t   � t e r s p e g l a   � n d r i n g a r   i   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g  V � r d :      A k t i v   s e s s i o n :   [ % d ]   % s  S e s s i o n   ' % s '   a v s l u t a d .  L o k a l   ' % s '   % s   F j � r r   ' % s '  ' % s '   b o r t t a g e n 7 � v e r v a k a r   f � r � n d r i n g a r ,   t r y c k   C T R L - C   f � r   a t t   a v b r y t a . . .  & H o p p a   � v e r   a l l a  K � r   g o d t y c k l i g t   f j � r r k o m m a n d o  & T e x t  & B i n � r t   8 � v e r f � r i n g s t y p :   % s | B i n � r | T e x t | A u t o m a t i s k   ( % s ) | A u t o m a t i s k O F i l n a m n s f � r � n d r i n g :   % s | I n g e n   � n d r i n g | V e r s a l e r | G e m e n e r | F � r s t a   v e r s a l | G e m e n e r   8 . 3  S � t t   r � t t i g h e t e r :   % s  L � g g   t i l l   X   t i l l   k a t a l o g  B e v a r a   t i d s s t � m p e l    F i l m a s k :   % s  R e n s a   ' A r k i v '   a t t r i b u t  B y t   i n t e   u t   o g i l t i g a   t e c k e n    B e v a r a   i n t e   t i d s s t � m p e l  B e r � k n a   i n t e   � v e r f � r i n g s s t o r l e k   S t a n d a r d � v e r f � r i n g s i n s t � l l n i n g a r  V � r d n a m n :   % s  A n v � n d a r n a m n :   % s  F j � r r k a t a l o g :   % s    L o k a l   k a t a l o g :   % s $ S k a n n a r   ' % s '   e f t e r   u n d e r k a t a l o g e r . . . % � v e r v a k a r   � n d r i n g a r   i   % d   k a t a l o g e r . . .  � n d r i n g   i   ' % s '   u p p t � c k t .  F i l   ' % s '   � v e r f � r d .  F i l   ' % s '   b o r t t a g e n . U % s   k o n f i g u r e r a d   � v e r f � r i n g s i n s t � l l n i n g   k a n   i n t e   a n v � n d a s   i   a k t u e l l   k o n t e x t | N � g o n | A l l a    I g n o r e r a   r � t t i g h e t s f e l  A n v � n d e r   a n v � n d a r n a m n   " % s " . . A n v � n d e r   t a n g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s " .  F e l a k t i g   l � s e n o r d .  � t k o m s t   n e k a d . 0 A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s "   f r � n   a g e n t . ( F � r s � k e r   m e d   p u b l i k   n y c k e l a u t e n t i s e r i n g . ' A u t e n t i s e r i n g   m e d   f � r i n s t � l l t   l � s e n o r d .  � p p n a r   t u n n e l . . .  A n s l u t n i n g   a v s l u t a d .    S � k e r   e f t e r   v � r d . . .  A n s l u t e r   t i l l   v � r d . . .  A u t e n t i s e r a r . . .  A u t e n t i s e r a d .  S t a r t a r   s e s s i o n e n . . .  L � s e r   f j � r r k a t a l o g . . .  S e s s i o n e n   s t a r t a d .  A n s l u t e r   g e n o m   t u n n e l . . .  S e r v e r   n e k a r   v � r   n y c k e l .  A d m i n i s t r a t i v t   f � r b j u d e n   ( % s ) .  A n s l u t n i n g   m i s s l y c k a d e s   ( % s ) . . N � t v e r k s f e l :   A n s l u t n i n g   t i l l   " % H O S T % "   n e k a d e s .   + N � t v e r k s f e l :   A n s l u t n i n g   � t e r s t � l l d   a v   p e e r . 5 N � t v e r k s f e l :   A n s l u t n i n g   t i l l   " % H O S T % "   g j o r d e   t i m e o u t . 2 V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s 
 & � t e r u p p t a / S e r v e r n   s t � d e r   i n t e   n � g r a   e x t r a   F T P   e g e n s k a p e r . . S e r v e r n   s t � d e r   d e   h � r   e x t r a   F T P   e g e n s k a p e r n a :   # � v e r f � r i n g s h a s t i g h e t s g r � n s :   % u   k B / s  & K o p i e r a   n y c k e l 
 & U p p d a t e r a 
 & L � g g   t i l l  B e v a r a   e n d a s t   l � s n i n g 	 J � m f � r . . .  S y n k r o n i s e r a r . . .  I n g e t   a t t   s y n k r o n i s e r a . 
 O b e g r � n s a d  S S L / T L S   I m p l i c i t   k r y p t e r i n g      T L S / S S L   E x p l i c i t   k r y p t e r i n g  V i s a r   a r g u m e n t e n   s o m   m e d d e l a n d e  H � m t a r   a t t r i b u t   f � r   f j � r r f i l # V � r d e n s   f i n g e r a v t r y c k s n y c k e l   � r   % s . F V � x e l   - f i l e m a s k   � s i d o s � t t e r   f � r � l d r a d e   i n k l u d e r a / e x k l u d e r a   a l t e r n a t i v .  B a r a   & n y a   o c h   � n d r a d e   f i l e r � S e r v e r n   a v v i s a d e   S F T P - a n s l u t n i n g ,   m e n   d e n   l y s s n a r   p �   F T P - a n s l u t n i n g a r . 
 
 V i l l   d u   a n v � n d a   F T P - p r o t o k o l l e t   i s t � l l e t   f � r   S F T P ?   F � r e d r a r   a t t   a n v � n d a   k r y p t e r i n g . ` � p p n a   s e s s i o n   m e d   k o m m a n d o r a d s p a r a m e t e r   i   s k r i p t   � r   f � r � l d r a d .   A n v � n d   ' o p e n ' - k o m m a n d o t   i s t � l l e t . L V A R N I N G !   A t t   g e   u p p   s � k e r h e t e n   o c h   a c c e p t e r a   n � g o n   n y c k e l   s o m   k o n f i g u r e r a t s ! P V A R N I N G !   A t t   g e   u p p   s � k e r h e t e n   o c h   a c c e p t e r a   n � g o t   c e r t i f i k a t   s o m   k o n f i g u r e r a t s !  N y   l o k a l   f i l   % s  N y   f j � r r f i l   % s $ L o k a l   f i l   % s   � r   n y a r e   � r   f j � r r f i l   % s $ F j � r r f i l   % s   � r   n y a r e   � n   l o k a l   f i l   % s  � v e r g e   f j � r r f i l   % s  � v e r g e   l o k a l   f i l   % s  S k i l l n a d e r   h i t t a d e :  T a   b o r t   E O F - t e c k e n  T a   b o r t   B O M [ A n v � n d a   k o n f i g u r e r a d e   � v e r f � r i n g s i n s t � l l n i n g a r   s o m   s k i l j e r   s i g   f r � n   f a b r i k s i n s t � l l n i n g a r n a . \ A n v � n d a   k o n f i g u r e r a d e   s y n k r o n i s e r i n g s a l t e r n a t i v   s o m   s k i l j e r   s i g   f r � n   f a b r i k s i n s t � l l n i n g a r n a .    V e r s i o n  U t v e c k l i n g s v e r s i o n  F e l s � k n i n g s v e r s i o n  -   D i s t r i b u e r a   I N T E ' S e r v e r n   s t � d e r   d e s s a   W e b D A V   u t � k n i n g a r :  E x k l u d e r a   & k a t a l o g e r " B e r � k n a r   k o n t r o l l s u m m a   a v   f j � r r f i l    L a d d a r   k l i e n t c e r t i f i k a t . . . < S e r v e r n   f r � g a r   e f t e r   a u t e n t i s e r i n g   m e d   e t t   k l i e n t c e r t i f i k a t .  L � s t  K � r b a r � S k r i p t   a n v � n d e r   i n t e   f r i s t � e n d e   p a r a m e t r a r .   P a r a m e t r a r n a   d u   h a r   a n g e t t   p �   k o m m a n d o r a d e n   k o m m e r   i n t e   a t t   a n v � n d a s .   D i n   k o m m a n d o r a d s y n t a x   � r   f � r m o d l i g e n   f e l . Z I   s k r i p t ,   b � r   d u   a n v � n d a   e n   - h o s t k e y   v � x e l   f � r   a t t   k o n f i g u r e r a   d e n   f � r v � n t a d e   v � r d n y c k e l n . Y I   s k r i p t   s k a   d u   i n t e   f � r l i t a   d i g   p �   s p a r a d e   w e b b p l a t s e r ,   a n v � n d a   d e t t a   k o m m a n d o   i s t � l l e t :  K o n f i g u r e r a   s e s s i o n s a l t e r n a t i v  A n s l u t    L a d d a   W i n S C P   . N E T   a s s e m b l e r  % s   ( i n k l u s i v e   k a t a l o g e r ) , F i l e n   m � s t e   v a r a   k o d a d   i   U T F - 8   e l l e r   U T F - 1 6 . 	 % s   o c h   % s  � n d r a r   l � s e n o r d .  & K l i s t r a   i n   n y c k e l  D u p l i c e r a r   f j � r r f i l e n    O k � n d ,         A l g o r i t m : 	 % s 
         S H A - 2 5 6 : 	 % s 
         M D 5 : 	 % s ) & K o p i e r a   n y c k e l f i n g e r a v t r y c k   t i l l   u r k l i p p . & K o p i e r a   c e r t i f i k a t   f i n g e r a v t r y c k   t i l l   u r k l i p p  K r y p t e r a   i n t e   n y a   f i l e r  E x k l u d e r a   d o l d a   f i l e r  E x k l u d e r a   t o m m a   k a t a l o g e r                                      C O R E _ V A R I A B L E ( S S H   o c h   S C P   k o d e n   � r   b a s e r a d   p �   P u T T Y   % s   " C o p y r i g h t   �   1 9 9 7  2 0 2 1   S i m o n   T a t h a m 3 h t t p s : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y /  F T P - k o d   b a s e r a d   p �   F i l e Z i l l a    C o p y r i g h t   �   T i m   K o s s e    h t t p s : / / f i l e z i l l a - p r o j e c t . o r g / m D e n n a   p r o d u k t   i n n e h � l l e r   p r o g r a m v a r a   s o m   u t v e c k l a t s   a v   O p e n S S L   P r o j e c t   f � r   a n v � n d n i n g   i   O p e n S S L : s   v e r k t y g   % s . ' C o p y r i g h t   �   1 9 9 8  % s   T h e   O p e n S S L   P r o j e c t    h t t p s : / / w w w . o p e n s s l . o r g / + W e b D A V / H T T P - k o d   b a s e r a d   p �   n e o n b i b l i o t e k   % s  C o p y r i g h t   �   1 9 9 9  2 0 2 0   J o e   O r t o n  h t t p s : / / n o t r o j . g i t h u b . i o / n e o n /  e X p a t   l i b r a r y   % s    h t t p s : / / l i b e x p a t . g i t h u b . i o /               ? h t t p s : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y / l i c e n c e . h t m l            * *  $ $ $ S 3 - k o d   b a s e r a d   p �   l i b s 3 - b i b l i o t e k   % s  C o p y r i g h t   �   B r y a n   I s c h o  h t t p s : / / g i t h u b . c o m / b j i / l i b s 3 0 h t t p s : / / g i t h u b . c o m / b j i / l i b s 3 / b l o b / m a s t e r / L I C E N S E                               & F e l   v i d   h � m t n i n g   a v   f i l l i s t a   f � r   " % s " . g C e r t i f i k a t   u t f � r d a d e s   i n t e   f � r   d e n   h � r   s e r v e r n .   D u   k a n s k e   a n s l u t e r   t i l l   e n   s e r v e r   s o m   l � t s a s   v a r a   " % s " . " I n g e n   f i l   m a t c h a n d e   ' % s '   h i t t a d e s . 0 V i s s a   c e r t i f i k a t   i   c e r t i f i k a t k e d j a n   � r   o g i l t i g a .    C e r t i f i k a t e t   � r   g i l t i g t . ! W e b D A V - r e s u r s   f l y t t a d e   t i l l   ' % s ' .  F � r   m � n g a   o m d i r i g e r i n g a r .  O m d i r i g e r i n g s l o o p   u p p t � c k t .  O g i l t i g   U R L   " % s " . ! P r o x y - a u t e n t i s e r i n g   m i s s l y c k a d e s . 1 V � r d n y c k e l   m a t c h a r   i n t e   k o n f i g u r e r a d   n y c k e l   " % s " ! < D e t   a n g i v n a   n a m n e t   k a n   i n t e   t i l l d e l a s   s o m   � g a r e   t i l l   e n   f i l . I D e t   a n g i v n a   n a m n e t   k a n   i n t e   t i l l d e l a s   s o m   d e n   p r i m � r a   g r u p p e n   f � r   e n   f i l . g D e n   b e g � r d a   � t g � r d e n   k u n d e   i n t e   s l u t f � r a s   e f t e r s o m   d e t   a n g i v n a   b y t e - i n t e r v a l l s l � s e t   i n t e   h a r   b e v i l j a t s . 7 P r i v a t   n y c k e l f i l   ' % s '   f i n n s   i n t e   e l l e r   k a n   i n t e   � p p n a s . & K o n t r o l l s u m m s a l g o r i t m   ' % s '   s t � d s   i n t e .  % s   % s   h a r   i n t e   v e r i f i e r a t s !   V a n l i g a   o r s a k e r   f � r   F e l k o d   4   � r : 
 -   B y t a   n a m n   p �   e n   f i l   t i l l   e t t   r e d a n   e x i s t e r a n d e   n a m n . 
 -   S k a p a   e n   k a t a l o g   s o m   r e d a n   f i n n s . 
 -   F l y t t a   e n   f j � r r f i l   t i l l   e t t   a n n a t   f i l s y s t e m   ( H D D ) . 
 -   � v e r f � r a   e n   f i l   t i l l   e t t   f u l l s t � n d i g t   f i l s y s t e m   ( H D D ) . 
 -   � v e r s k r i d a   e n   a n v � n d a r e s   d i s k k v o t .  K a n   i n t e   � p p n a   c e r t i f i k a t   " % s " .    K a n   i n t e   l � s a   c e r t i f i k a t   " % s " .   F e l   v i d   a v k o d n i n g   a v   c e r t i f i k a t . % F e l   v i d   a v k o d n i n g   a v   c e r t i f i k a t   " % s " . c C e r t i f i k a t f i l e n   " % s "   i n n e h � l l e r   i n t e   e n   p u b l i k   n y c k e l   o c h   i n g e n   m o t s v a r a n d e   . c r t / . c e r - f i l   h i t t a d e s .  F e l   v i d   l � s n i n g   a v   f i l e n   ' % s ' . ! F e l   v i d   u p p l � s n i n g   a v   f i l e n   ' % s ' .  F i l e n   ' % s '   � r   i n t e   l � s t . ) F e l   v i d   s p a r a n d e   a v   n y c k e l   t i l l   f i l   " % s " . K N e o n   H T T P - b i b l i o t e k e t s   i n i t i a l i s e r i n g   m i s s l y c k a d e s ,   k a n   i n t e   � p p n a   s e s s i o n . � V � l j a   f i l e r   m e d   h j � l p   a v   e t t   s � k v � g s s l u t   m e d   s n e d s t r e c k   � r   t v e t y d i g .   T a   b o r t   s n e d s t r e c k e t   f � r   a t t   v � l j a   m a p p .   B i f o g a   *   m a s k   f � r   a t t   v � l j a   a l l a   f i l e r   i   m a p p e n . � N � r   d u   a n s l u t e r   m e d   h j � l p   a v   e n   I P - a d r e s s ,   � r   d e t   i n t e   m � j l i g t   a t t   k o n t r o l l e r a   o m   c e r t i f i k a t e t   u t f � r d a d e s   f � r   s e r v e r n .   A n v � n d   e t t   v � r d n a m n   i s t � l l e t   f � r   I P - a d r e s s e n . E F � r v � n t a d e   v � r d n y c k e l   h a r   i n t e   k o n f i g u r e r a t s ,   a n v � n d   - h o s t k e y   s w i t c h . * O m d i r i g e r a s   t i l l   e n   o k r y p t e r a d   w e b b a d r e s s .  M o t t o g   s v a r   % d   " % s "   f r � n   % s . 2 F i l e Z i l l a   w e b b p l a t s h a n t e r a r f i l   h i t t a d e s   i n t e   ( % s ) . @ I n g a   w e b b p l a t s e r   h i t t a d e s   i   F i l e Z i l l a   w e b b p l a t s h a n t e r a r f i l   ( % s ) . ' F i l e Z i l l a   w e b b p l a t s   " % s "   h i t t a d e s   i n t e . [ D u   k a n   i n t e   a n s l u t a   t i l l   e n   S F T P - s e r v e r   m e d   h j � l p   a v   e n   F T P - p r o t o k o l l .   V � l j   r � t t   p r o t o k o l l . - F e l   u p p s t o d   v i d   l o g g n i n g .   K a n   i n t e   f o r t s � t t a .  ' % s '   � r   i n t e   e n   g i l t i g   s t o r l e k . ( O p e n S S H   f i l e n   k n o w n _ h o s t s   h i t t a d e s   i n t e . % I n g a   v � r d n y c k l a r   f i n n s   i   k n o w n _ h o s t s . R U r k l i p p e t s   i n n e h � l l   s t � m m e r   i n t e   � v e r e n s   m e d   v � r d n y c k e l n   e l l e r   d e s s   f i n g e r a v t r y c k . 
 R e s u r s :   % s  Y t t e r l i g a r e   d e t a l j e r :   % s  E x t r a   d e t a l j e r :  � t k o m s t   n e k a d . / F i l e n   � r   i n t e   k r y p t e r a d   m e d   e n   k � n d   k r y p t e r i n g . � * * O g i l t i g   k r y p t e r i n g s n y c k e l . * * 
 
 K r y p t e r i n g s n y c k e l n   f � r   k r y p t e r i n g   % s   m � s t e   h a   % d   b y t e .   D e n   m � s t e   a n g e s   i   h e x a d e c i m a l   r e p r e s e n t a t i o n   ( d v s   % d   t e c k e n ) . ) S e r v e r   s k i c k a d e   e n   f i l   s o m   i n t e   b e g � r d e s . & D e t   g i c k   i n t e   a t t   l a g r a   n y   v � r d n y c k e l . [ N � r   d u   l a d d a r   u p p   s t r e a m a d   d a t a   k a n   e n d a s t   e n   k � l l a   a n g e s   o c h   m � l e t   m � s t e   a n g e   e t t   f i l n a m n .   # F e l   v i d   l � s n i n g   a v   i n m a t n i n g s s t r � m .                                                         	 W I N _ E R R O R   Q % s 
   
 V a r n i n g :   A t t   a v b r y t a   d e n   h � r   o p e r a t i o n e n   k o m m e r   a t t   s t � n g a   n e r   a n s l u t n i n g e n !          K a n   i n t e   s k a p a   g e n v � g . ) K a n   i n t e   s k r i v a   � v e r   s p e c i a l s e s s i o n   ' % s ' .  K a n   i n t e   u t f o r s k a   k a t a l o g   ' % s ' . + I n g e n   f i l l i s t a   f � r   � v e r f � r i n g   h a r   a n g i v i t s .  K a n   i n t e   s k a p a   k a t a l o g e n   ' % s ' .   ' K a n   i n t e   t a   b o r t   t e m p o r � r   k a t a l o g   ' % s ' . % K a n   i n t e   � p p n a   e l l e r   k � r a   f i l e n   ' % s ' .  K a n   i n t e   s t a r t a   e d i t o r   ' % s ' .   w K a n   i n t e   � p p n a   m o t s v a r a d e   k a t a l o g   i   m o t s a t t   p a n e l .   S y n k r o n i s e r i n g   a v   k a t a l o g b l � d d r i n g   m i s s l y c k a d e s .   D e n   h a r   s t � n g t s   a v .  K a n   i n t e   a v g � r a   g e n v � g   ' % s ' .   % ' % s '   � r   i n t e   g i l t i g t   p r o f i l p l a t s n a m n . 4 ' % s '   � r   i n t e   g i l t i g t   n a m n   f � r   e n   p r o f i l p l a t s k a t a l o g . 1 P r o f i l p l a t s k a t a l o g e n   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . 5 B e s k r i v n i n g   p �   e g e t   k o m m a n d o   k a n   i n t e   i n n e h � l l a   ' % s ' . 1 E g e t   k o m m a n d o   m e d   b e s k r i v n i n g e n   ' % s '   f i n n s   r e d a n . D K a n   i n t e   f r � g a   a p p l i k a t i o n e n s   h e m s i d a   e f t e r   u p p d a t e r i n g s i n f o r m a t i o n . , F e l   u p p s t o d   v i d   s � k n i n g   e f t e r   u p p d a t e r i n g a r .         < K a n   i n t e   r e g i s t r e r a   p r o g r a m m e t   f � r   a t t   h a n t e r a   U R L - a d r e s s e r . 2 M u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . E S k a l   d r a - t i l l � g g e t   m u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . �* * W i n S C P   k u n d e   i n t e   i d e n t i f i e r a   k a t a l o g e n ,   s o m   f i l e n   s l � p p t e s   i . * *   A n t i n g e n   h a r   d u   i n t e   s l � p p t   f i l e n   i   e n   v a n l i g   k a t a l o g   ( t . e x .   U t f o r s k a r e n )   e l l e r   o m   d u   i n t e   h a r   s t a r t a t   o m   d a t o r n   � n n u   e f t e r   i n s t a l l a t i o n e n   a v   s k a l t i l l � g g e t   d r a   &   s l � p p .   
 
 A l t e r n a t i v t   k a n   d u   v � x l a   t i l l   k o m p a t i b e l   d r a   &   s l � p p l � g e   ( f r � n   i n s t � l l n i n g s f � n s t r e t ) ,   s o m   a n v � n d e r   t e m p o r � r a   k a t a l o g e r   f � r   n e d l a d d n i n g a r .   D e t   g � r   a t t   d u   s l � p p a   f i l e r   t i l l   a l l a   d e s t i n a t i o n e r . K F i l e n   ' % s '   i n n e h � l l e r   i n t e   n � g o n   � v e r s � t t n i n g   f � r   d e n   h � r   p r o d u k t v e r s i o n e n . 5 F i l e n   ' % s '   i n n e h � l l e r   � v e r s � t t n i n g   f � r   % s   v e r s i o n   % s .   8 G S S A P I / S S P I   m e d   K e r b e r o s   s t � d s   i n t e   p �   d e t   h � r   s y s t e m e t . ' F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r . 8 F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r   i   k a t a l o g e n   ' % s ' .   6 F e l   u p p s t o d   v i d   b e v a k n i n g e n   a v   � n d r i n g a r   i   f i l e n   ' % s ' . � * * K a n   i n t e   � v e r f � r a   d e n   r e d i g e r a d e   f i l e n   ' % s ' * * 
 
 S e s s i o n e n   ' % s '   h a r   r e d a n   s t � n g t s . 
 
 � p p n a   e n   n y   s e s s i o n   p �   s a m m a   w e b b p l a t s   o c h   f � r s � k   s p a r a   f i l e n   i g e n . I D e t   f i n n s   r e d a n   f � r   m � n g a   f i l e r   � p p n a d e .   V a r   g o d   s t � n g   n � g r a   f i l e r   f � r s t .   R % s   V a r   v � n l i g   t a   b o r t   f i l e n .   A n n a r s   k o m m e r   i n t e   a p p l i k a t i o n e n   a t t   f u n g e r a   k o r r e k t . o K a n   i n t e   s k a p a   t e m p o r � r   k a t a l o g   ' % s ' .   D u   k a n   � n d r a   r o t k a t a l o g e n   f � r   l a g r i n g   a v   t e m p o r � r a   f i l e r   i   I n s t � l l n i n g a r . �W i n S C P   k u n d e   i n t e   a v g � r a   v i l k e t   p r o g r a m   s o m   s k a   s t a r t a s   f � r   a t t   � p p n a   f i l e n .   W i n S C P   k a n   i n t e   b e v a k a   � n d r i n g a r   i   f i l e n ,   s �   d e n   v i l l   i n t e   l a d d a s   u p p . 
   
 E n   m � j l i g   o r s a k   t i l l   p r o b l e m e t   � r   a t t   f i l e n   r e d a n   h a r   � p p n a t s   a v   e t t   a n n a t   p r o g r a m   s o m   k � r s . 
   
 O m   d u   v i l l   a n v � n d a   p r o g r a m m e t   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r . 
   
 N o t e r a   a t t   f i l e n   l i g g e r   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . � N � g r a   a v   d e   t e m p o r � r a   k a t a l o g e r n a   k u n d e   i n t e   t a s   b o r t .   O m   f i l e r   f i n n s   l a g r a d e   d � r   s o m   f o r t f a r a n d e   � r   � p p n a ,   s t � n g   d e s s a   o c h   p r o v a   i g e n . � F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o ,   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   e n a   p a n e l e n ,   f � r   a t t   k � r a   k o m m a n d o t   p �   d e   v a l d a   f i l e r n a   i   m o t s a t t   p a n e l .   A l t e r n a t i v t   k a n   s a m m a   a n t a l   f i l e r   m a r k e r a s   i   b � d a   p a n e l e r n a   f � r   a t t   k � r a   k o m m a n d o t   p �   m a t c h a n d e   p a r   a v   f i l e r . W F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o t   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   l o k a l a   p a n e l e n . � N � g r a   a v   d e   v a l d a   f j � r r f i l e r n a   l a d d a d e s   i n t e   n e r .   D e t   v a l d a   e g n a   k o m m a n d o t   m � s t e   k � r a s   p �   m a t c h a n d e   p a r   a v   f i l e r ,   v i l k e t   d � r f � r   i n t e   � r   m � j l i g t . $ K a n   i n t e   i n i t i a l i s e r a   e x t e r n   k o n s o l .   N K a n   i n t e   � p p n a   m a p p n i n g s o b j e k t   f � r   a t t   s t a r t a   k o m m u n i k a t i o n   m e d   e x t e r n   k o n s o l . ; T i m e o u t   v � n t a r   p �   e x t e r n   k o n s o l   f � r   a t t   s l u t f � r a   k o m m a n d o t . 4 I n k o m p a t i b e l t   p r o t o k o l l v e r s i o n   f � r   e x t e r n   k o n s o l   % d . D F e l   u p p s t o d   n � r   s � k v � g   ' % s '   l a d e s   t i l l   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) . H F e l   u p p s t o d   n � r   s � k v � g   ' % s '   t o g s   b o r t   f r � n   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) .   [ F i l e n   ' % s '   � r   r e d a n   � p p n a d   i   e n   e x t e r n   e d i t o r   ( a p p l i k a t i o n )   e l l e r   h � l l e r   p �   a t t   l a d d a s   u p p . 8 D u   h a r   i n t e   a n g i v i t   n � g o n   a u t o m a t i s k t   v a l   a v   m a s k r e g l e r . D F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   m e d   b e s k r i v n i n g   ' % s '   f i n n s   r e d a n . x * * A n p a s s a t   k o m m a n d o   ' % s '   k a n   i n t e   k � r a s   j u s t   n u . * *   D u   k a n   b e h � v a   v � l j a   f i l e r   f � r   k o m m a n d o t   e l l e r   � p p n a   e n   s e s s i o n   f � r s t . A K a n   i n t e   l a d d a   o m   f i l e n   ' % s ' ,   s e s s i o n e n   ' % s '   h a r   r e d a n   a v s l u t a t s .         L � s e n o r d e t   k a n   i n t e   d e k r y p t e r a s . 3 D u   h a r   i n t e   a n g e t t   k o r r e k t   n u v a r a n d e   h u v u d l � s e n o r d . 0 N y a   o c h   u p p r e p a d e   h u v u d l � s e n o r d e t   � r   i n t e   s a m m a .   F E x t e r n   k o n s o l u t d a t a   d i r i g e r a s   t i l l   p i p e .   S e   t i l l   a t t   p i p e n   l � s e s   f r � n . ) ' % s '   � r   a r b e t s y t a ,   i n t e   w e b b p l a t s k a t a l o g . ) ' % s '   � r   w e b b p l a t s k a t a l o g ,   i n t e   a r b e t s y t a . ) F e l   v i d   e x e k v e r i n g   a v   k o m m a n d o   " % s "   ( % s ) . A K a n   i n t e   l � g g a   t i l l   s � k v � g   t i l l   % P A T H % ,   % P A T H %   � r   r e d a n   f � r   l � n g . 
 S t a c k s p � r :     ? I n g a   w e b b p l a t s e r   h i t t a d e s   i   P u T T Y   w e b b p l a t s r e g i s t e r n y c k e l   ( % s ) .   I n g e n   w e b b p l a t s m a s k   s p e c i f i c e r a d * I n g a   w e b b p l a t s i n s t � l l n i n g a r   s p e c i f i c e r a d e .  I n t e   � n d r a d    � n d r a d . H i t t a d e   % d   w e b b p l a t s e r ,   � n d r a d e   % d   w e b b p l a t s e r ! D u   m � s t e   a n g e   i n g � e n d e   n y c k e l f i l .  I n g e n   � t g � r d   a n g i v e n . " R e d i g e r a   S S H - 1   n y c k l a r   s t � d s   i n t e .  L � s e n f r a s e r n a   m a t c h a r   i n t e . ! D u   m � s t e   a n g e   u t g � e n d e   n y c k e l f i l . 4 F e l   v i d   h � m t n i n g   a v   u p p d a t e r i n g .   F � r s � k   i g e n   s e n a r e . E D e n   n e d l a d d a d e   u p p d a t e r i n g   k u n d e   i n t e   v e r i f i e r a s .   F � r s � k   i g e n   s e n a r e . C D i n   e - p o s t a d r e s s   h a r   i n t e   b e h � r i g h e t   f � r   a u t o m a t i s k a   u p p d a t e r i n g a r . F D i n   e - p o s t a d r e s s   b e h � r i g h e t   f � r   a u t o m a t i s k a   u p p d a t e r i n g a r   h a r   u p p h � r t . ^ D i n   e - p o s t a d r e s s   b l o c k e r a d e s   t i l l   a u t o m a t i s k a   u p p d a t e r i n g a r   p �   g r u n d   a v   � v e r d r i v e n   a n v � n d n i n g . � F � r   a t t   a k t i v e r a   a u t o m a t i s k a   u p p d a t e r i n g a r   f � r   d i n   e - p o s t a d r e s s ,   v � n l i g e n   f y l l   i   e t t   d o n a t i o n s f o r m u l � r   ( i n k l u s i v e   d i n   p o s t a d r e s s ) . 
 
 D u   h i t t a r   e n   l � n k   t i l l   f o r m u l � r e t   i   e t t   k v i t t o   s o m   d u   h a r   f � t t   e f t e r   d i n   d o n a t i o n . U D i n   d o n a t i o n   � r   u n d e r   d e n   g r � n s   s o m   k r � v s   f � r   a t t   a k t i v e r a   a u t o m a t i s k a   u p p d a t e r i n g a r . 
 I n g a   t i p s . & K o n v e r t e r a   p u b l i k a   n y c k l a r   s t � d s   i n t e .   / S � k e r   s e s s i o n   ( S S H   e l l e r   T L S / S S L )   i n t e   a n g i v e n .  U t � k n i n g e n   k r � v e r   % s . / O g i l t i g t   v � r d e   " % s "   f � r   u t � k n i n g s d i r e k t i v e t   % s . * S a k n a r   o b l i g a t o r i s k t   u t � k n i n g s d i r e k t i v   % s . " I n g e n   u t � k n i n g   f i n n s   i   d o k u m e n t e t . , D e t   f i n n s   r e d a n   e n   u t � k n i n g   m e d   n a m n e t   " % s " .   U t � k n i n g e n   � r   r e d a n   i n s t a l l e r a d . + F e l   v i d   i n l � s n i n g   a v   e n   u t � k n i n g   f r � n   " % s " . i * * I n g e n   s e s s i o n   � r   � p p e n * * 
 D e t   v a l d a   k o m m a n d o t   h a r   p l a t s s p e c i f i k a   a l t e r n a t i v ,   m e n   i n g e n   s e s s i o n   � r   � p p e n . (* * W i n S C P   k u n d e   i n t e   u p p t � c k a   e n   m a p p   d � r   d e   s l � p p t a   f i l e r n a   s l � p p t e s . * *   I   s t a n d a r d l � g e t   f � r   D r a   o c h   s l � p p   t i l l � t e r   W i n S C P   a t t   e n d a s t   f i l e r   s l � p p s   t i l l   l o k a l a   e n h e t e r   o c h   m a p p a d e   n � t v e r k s e n h e t e r . 
 
 D u   k a n   t i l l � t a   a t t   f i l e r   s l � p p s   t i l l   a n d r a   m � l   i   i n s t � l l n i n g a r .   T r y c k   p �   H j � l p - k n a p p e n   f � r   d e t a l j e r . " F e l   v i d   u p p d a t e r i n g   a v   s n a b b l i s t a .                      W I N _ C O N F I R M A T I O N . S e s s i o n   m e d   n a m n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ! K a t a l o g e n   ' % s '   f i n n s   i n t e .   S k a p a ?   � * * A v b r y t   f i l � v e r f � r i n g ? * * 
   
 O p e r a t i o n e n   k a n   i n t e   a v b r y t a s   i   m i t t e n   a v   f i l � v e r f � r i n g . 
 T r y c k   ' J a '   f � r   a t t   a v b r y t a   f i l � v e r f � r i n g   o c h   s t � n g a   a n s l u t n i n g e n . 
 T r y c k   ' N e j '   F � r   a t t   a v s l u t a   a k t u e l l   f i l � v e r f � r i n g . 
 T r y c k   ' A v b r y t '   f � r   a t t   f o r t s � t t a   o p e r a t i o n e n . . � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   f i l e n   ' % s ' ? 7 � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   d e   % d   v a l d a   f i l e r n a ? / A v s l u t a   s e s s i o n e n   ' % s '   o c h   s t � n g   a p p l i k a t i o n e n ?  F r � g a   m i & g   a l d r i g   i g e n 9F � r   l i t e   l e d i g t   u t r y m m e   p �   t e m p o r � r   e n h e t ! 
 
 N � r   f i l e r   d r a s   f r � n   e n   f j � r r k a t a l o g ,   l a d d a s   f i l e r n a   f � r s t   n e r   t i l l   e n   t e m p o r � r   k a t a l o g   ' % s ' .   D e t   � r   % s   l e d i g t   p �   e n h e t e n .   T o t a l   s t o r l e k   f � r   d e   v a l d a   f i l e r n a   � r   % s . 
 
 O B S :   T e m p o r � r   k a t a l o g e n   k a n   � n d r a s   i   I n s t � l l n i n g s f � n s t r e t . 
 
 V i l l   d u   f o r t s � t t a   m e d   a t t   l a d d a   n e r   f i l e r n a ?   ( L � g g   t i l l   k a t a l o g e n   ' % s '   t i l l   b o k m � r k e n ?     - S k a p a   g e n v � g   p �   s k r i v b o r d e t   f � r   s e s s i o n   ' % s ' ? 2 A n v � n d   a k t u e l l a   s e s s i o n s i n t � l l n i n g a r   s o m   s t a n d a r d ?  & H o p p a   � v e r # F i l e n   h a r   � n d r a t s .   S p a r a   � n d r i n g a r ? 9 S k a p a   u t f o r s k a r e n s   ' S k i c k a   t i l l ' - g e n v � g   f � r   s e s s i o n   ' % s ' ?  S k a p a   v a l d   i k o n / g e n v � g ? / A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   a p p l i k a t i o n e n ?   T a   b o r t   v a l d   p r o f i l p l a t s k a t a l o g ?  & F � r e g � e n d e  & N � s t a   3 V i l l   d u   r e g i s t r e r a   W i n S C P   a t t   h a n t e r a   U R L - a d r e s s e r ? L V i l l   d u   r e n s a   u p p   d a t a   f r � n   d e n   h � r   d a t o r n   s o m   h a r   s k a p a t s   a v   a p p l i k a t i o n e n ? ! % s 
 
 V i l l   d u   s t � n g a   a p p l i k a t i o n e n ? G % % s 
 
 V i l l   d u   a v s l u t a   % d   � t e r s t � e n d e   s e s s i o n e r   o c h   s t � n g a   a p p l i k a t i o n e n ? � * * D e t   f i n n s   f o r t f a r a n d e   n � g r a   � v e r f � r i n g a r   i   b a k g r u n d s k � n .   V i l l   d u   k o p p l a   n e r   i a l l a f a l l ? * * 
 
 V a r n i n g :   O m   d u   t r y c k e r   p �   ' O K '   k o m m e r   a l l a   � v e r f � r i n g a r   a t t   a v s l u t a s   o m e d e l b a r t . * * V i l l   d u   � p p n a   s e p a r a t   s k a l s e s s i o n ? * * 
 
 N u v a r a n d e   s e s s i o n   % s   s t � d e r   i n t e   k o m m a n d o t   d u   b e g � r .   S e p a r a t   s k a l s e s s i o n   k a n   � p p n a s   f � r   a t t   b e a r b e t a   k o m m a n d o t . 
 
 O B S :   S e r v e r n   m � s t e   e r b j u d a   U n i x - l i k n a n d e   s k a l   o c h   s k a l e t   m � s t e   a n v � n d a   s a m m a   s � k v � g s s y n t a x   s o m   n u v a r a n d e   s e s s i o n   % s . � D e t   f i n n s   n � g r a   � p p n a   f i l e r .   V a r   v � n l i g   s t � n g   d e m   i n n a n   a p p l i k a t i o n e n   a v s l u t a s . 
   
 O B S :   O m   d e t t a   i n t e   u t f � r s ,   k a n   r e d i g e r a d e   f i l e r   l i g g a   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . '* * V i l l   d u   t a   b o r t   t i d i g a r e   t i l l f � l l i g a   k a t a l o g e r ? * * 
 
 W i n S C P   h a r   h i t t a t   % d   t e m p o r � r a   k a t a l o g e r ,   s o m   f � r m o d l i g e n   h a r   s k a p a t s   t i d i g a r e .   D e s s a   k a t a l o g e r   k a n   i n n e h � l l a   f i l e r   s o m   t i d i g a r e   h a r   r e d i g e r a t s   e l l e r   l a d d a t s   n e r . 
 
 D u   k a n   o c k s �   � p p n a   k a t a l o g e r   f � r   a t t   s e   � v e r   i n n e h � l l e t   o c h   t a   b o r t   d e m   s j � l v .  & � p p n a # V i s a   i n t e   d e t   h � r   m e d d e l a n d e t   i & g e n   f * * V i l l   d u   s k a p a   s k r i v b o r d s i k o n   f � r   a l l a   a n v � n d a r e ? * * 
 
 D u   m � s t e   h a   a d m i n i s t r a t � r s r � t t i g h e t e r   f � r   d e t t a . U V i l l   d u   l � g g a   t i l l   a p p l i k a t i o n e n s   s � k v � g   ' % s '   t i l l   m i l j � v a r i a b e l n s   s � k v � g   ( % % P A T H % % ) ? �E d i t o r n   ( a p p l i k a t i o n )   s o m   s t a r t a d e s   f � r   a t t   � p p n a   f i l   ' % s '   a v s l u t a d e s   f � r   t i d i g t .   O m   d e n   i n t e   a v s l u t a d e s   a v   e r ,   k a n   d e t   b e r o   p �   a t t   d e n   e x t e r n a   e d i t o r   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   e d i t o r n   s k i c k a r   s e d a n   d e n   n y a   f i l e n   t i l l   b e f i n t l i g a   i n s t a n s e r   a v   e d i t o r n   o c h   a v s l u t a r   s i g   o m e d e l b a r t .   F � r   a t t   s t � d j a   d e n n a   t y p   a v   e d i t o r s ,   m � s t e   W i n S C P   a n p a s s a   s i t t   b e t e e n d e ,   i n t e   t a   b o r t   t e m p o r � r   f i l   n � r   p r o c e s s e n   a v s l u t a r ,   u t a n   a t t   b e h � l l a   d e n   s �   l � n g e   W i n S C P   � r   i g � n g .   B e t e e n d e t   k a n   s t � n g a s   a v   g e n o m   a t t   � n d r a   i n s t � l l n i n g a r   f � r   e d i t o r n   ' E x t e r n   e d i t o r   � p p n a r   v a r j e   f i l   i   e t t   s e p a r a t   f � n s t e r   ( p r o c e s s ) ' .   O m   d i n   e d i t o r   i n t e   � r   a v   d e t   h � r   s l a g e t ,   b o r t s e   f r � n   d e t t a   m e d d e l a n d e   o c h   l � t   f i l e n   t a s   b o r t   f r � n   d e n   t e m p o r � r a   k a t a l o g e n   n u . 
   
 V i l l   n i   t a   b o r t   d e n   � p p n a d e   f i l e n   n u ?   ( G e n o m   a t t   t r y c k a   p �   ' N e j '   k o m m e r   d u   a t t   m � j l i g g � r a   d e t   s � r s k i l d a   b e t e e n d e t   o c h   b e h � l l a   f i l e n   i   t e m p o r � r a   k a t a l o g e n . )   � * * V i l l   d u   g � r a   r i k t n i n g e n   d u   v a l t   t i l l   s t a n d a r d ? * * 
 
 D u   h a r   � s i d o s a t t   f � r v a l d   s y n k r o n i s e r i n g s r i k t n i n g .   S o m   s t a n d a r d   b e s t � m s   r i k t n i n g e n   a v   f i l p a n e l e n   s o m   v a r   a k t i v   i n n a n   i n n a n   d u   k � r d e   s y n k r o n i s e r i n g s f u n k t i o n e n . � * * V i l l   d u   f � r s t   u t f � r a   e n   f u l l s t � n d i g   s y n k r o n i s e r i n g   a v   f j � r r k a t a l o g e n ? * * 
 
 F u n k t i o n e n   ' H � l l   f j � r r k a t a l o g   u p p d a t e r a d '   f u n g e r a r   k o r r e k t   e n d a s t   o m   f j � r r k a t a l o g e n   � r   s y n k r o n i s e r a d   m e d   d e n   l o k a l a   i n n a n   d e n   s t a r t a r . 1 S � k e r   p �   a t t   d u   v i l l   t a   b o r t   s p a r a d   s e s s i o n   ' % s ' ? � F l e r   � n   % d   k a t a l o g e r   o c h   u n d e r k a t a l o g e r   h i t t a d e s .   B e v a k n i n g   a v   � n d r i n g a r   i   m � n g a   k a t a l o g e r   k a n   s i g n i f i k a n t   m i n s k a   p r e s t a n d a n   p �   d a t o r n . 
   
 V i l l   d u   s k a n n a   f l e r   k a t a l o g e r ,   u p p   t i l l   % d   k a t a l o g e r ? 	 % s   ( % d   s )   8 S � k e r   p �   a t t   d u   v i l l   f l y t t a   f i l   ' % s '   t i l l   p a p p e r s k o r g e n ? > S � k e r   p �   a t t   d u   v i l l   f l y t t a   % d   v a l d a   f i l e r   t i l l   p a p p e r s k o r g e n ? I F i l e n   h a r   � n d r a t s .   � n d r i n g a r   v i l l   f � r l o r a s ,   o m   f i l e n   l a d d a s   o m .   F o r t s � t t ?  K & o n f i g u r e r a . . . ^ * * V i l l   d u   f � r s � k a   s k a p a   k a t a l o g e n   ' % s ' ? * * 
 
 K a n   i n t e   � p p n a   m o t s v a r a n d e   k a t a l o g   i   m o t s a t t   p a n e l .  L � g g   t i l l   & d e l a d e   b o k m � r k e n s* * V i l l   d u   s k i c k a   m e d d e l a n d e t   t i l l   W i n S C P : s   w e b b p l a t s ? * * 
 
 D e t   f i n n s   i n g e n   h j � l p s i d a   a s s o c i e r a d   m e d   m e d d e l a n d e t .   W i n S C P   k a n   s � k a   p �   s i n   d o k u m e n t a t i o n s p l a t s   e f t e r   m e d d e l a n d e t e x t e n . 
 
 O B S :   W i n S C P   k o m m e r   a t t   s k i c k a   m e d d e l a n d e t   � v e r   e n   o s � k e r   a n s l u t n i n g .   K o n t r o l l e r a   a t t   m e d d e l a n d e t   i n t e   i n n e h � l l e r   n � g o n   d a t a   s o m   d u   v i l l   s k y d d a ,   t i l l   e x e m p e l   n a m n   p �   f i l e r ,   k o n t o n   e l l e r   v � r d a r . 9* * D i t t   l � s e n o r d   � r   f � r   e n k e l t   o c h   k a n   i n t e   g e   t i l l r � c k l i g t   s k y d d   m o t   a t t a c k e r   m e d   o r d l i s t a   e l l e r   b r u t e   f o r c e . 
 � r   d u   s � k e r   a t t   d u   v i l l   a n v � n d a   d e t ? * * 
 
 O B S :   b r a   l � s e n o r d   h a r   m i n s t   s e x   t e c k e n   o c h   i n n e h � l l e r   b � d e   g e m e n e r   o c h   v e r s a l e r ,   s i f f r o r   o c h   s p e c i a l t e c k e n ,   s �   s o m   a v g r � n s a r e ,   s y m b o l e r ,   b o k s t � v e r   m e d   a c c e n t ,   e t c . 9 S k a p a   g e n v � g   p �   s k r i v b o r d e t   t i l l   w e b b p l a t s k a t a l o g e n   ' % s ' ? 0 S k a p a   g e n v � g   p �   s k r i v b o r d e t   t i l l   a r b e t s y t a   ' % s ' ? E V i l l   d u   � t e r a n s l u t a   s e s s i o n   ' % s '   f � r   a t t   � v e r f � r a   r e d i g e r a d   f i l   ' % s ' ? K A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   a p p l i k a t i o n e n   u t a n   a t t   s p a r a   e n   a r b e t s y t a ? � * * V i l l   d u   a n v � n d a   % s   i s t � l l e t   f � r   i n t e r n a   s t a n d a r d e d i t o r ? * * 
 
 W i n S C P   h a r   u p p t � c k t   a t t   d u   h a r   d e n   a n p a s s a d e   t e x t e d i t o r n   ' % s '   a s s o c i e r a d   m e d   t e x t f i l e r . � * * D u   h a r   s p a r a t   s e s s i o n e r / w e b b p l a t s e r   i   % s . 
 
 V i l l   d u   i m p o r t e r a   d e m   t i l l   W i n S C P ? * * 
 
 ( D u   k a n   i m p o r t e r a   d e m   n � r   s o m   h e l s t   s e n a r e   i   d i a l o g r u t a n   L o g g a   i n ) | P u T T Y   S S h - k l i e n t | F i l e z i l l a   F T P - k l i e n t | % s   o c h   % s k I m p o r t e r a   k o n f i g u r a t i o n   k o m m e r   a t t   s k r i v a   � v e r   a l l a   d i n a   i n s t � l l n i n g a r   o c h   w e b b p l a t s e r . 
 
 V i l l   d u   f o r t s � t t a ?  & A l l a    J & a   t i l l   a l l a  R a & p p o r t e r a � D e t   f i n n s   a n d r a   i n s t a n s e r   a v   W i n S C P   i g � n g . 
 
 S t � l l a   i n   e l l e r   r e n s a   h u v u d l � s e n o r d e t ,   m e d a n   e n   a n n a n   i n s t a n s   a v   W i n S C P   � r   i g � n g ,   k a n   o r s a k a   f � r l u s t   a v   d i n a   l a g r a d e   l � s e n o r d . 
 
 V � n l i g e n   a v s l u t a   a n d r a   i n s t a n s e r   a v   W i n S C P   i n n a n   d u   f o r t s � t t e r . � V i l l   d u   b i f o g a   r e d i g e r a d   f i l   ' % s '   t i l l   s e s s i o n   ' % s ' ? * * 
 
 O r i g i n a l   s e s s i o n e n   s o m   a n v � n d e s   f � r   a t t   l a d d a   n e r   f i l e n   ' % s '   t i l l   e d i t o r n   h a r   r e d a n   s t � n g t s . @ V i l l   d u   a v r e g i s t r e r a   W i n S C P   f r � n   h a n t e r i n g   a v   a l l a   U R L - a d r e s s e r ? * * F � r s � k   a t t   � p p n a   s t o r   f i l ? * * 
 
 F i l e n   d u   f � r s � k e r   � p p n a   i   e n   i n t e r n   e d i t o r   � r   f � r   s t o r   ( % s ) .   W i n S C P   i n t e r n   e d i t o r   � r   i n t e   a v s e d d   f � r   r e d i g e r i n g   a v   s t o r a   f i l e r .   � v e r v � g   a t t   a n v � n d a   e n   e x t e r n   e d i t o r   s o m   k a n   r e d i g e r a   s t o r a   f i l e r . 
 
 D u   k a n   f � r s � k a   � p p n a   f i l e n   � n d � ,   m e n   W i n S C P   k a n   m i s s l y c k a s .  S t � n g X U t � k n i n g e n   k o m m e r   i n t e   f r � n   e n   b e t r o d d   k � l l a .   � r   d u   s � k e r   p �   a t t   d u   v i l l   i n s t a l l e r a   d e n ? � * * A n v � n d e r   d e n   s e n a s t e   k o m p a t i b l a   o c h   b e t r o d d a   v e r s i o n   a v   u t � k n i n g e n . * * 
 
 D e n   s e n a s t e   v e r s i o n e n   a v   u t � k n i n g e n   h a r   a n t i n g e n   i n t e   g r a n s k a t s   e l l e r   � r   i n t e   k o m p a t i b e l   m e d   d e n   h � r   v e r s i o n e n   a v   W i n S C P . [* * V i l l   d u   s k r i v a   � v e r   e n   b e f i n t l i g   I N I - f i l   ' % s ' ? * * 
 
 V � l j   ' S k r i v   � v e r '   f � r   a t t   s k r i v a   � v e r   d e n   v a l d a   I N I - f i l e n   m e d   d e n   a k t u e l l a   k o n f i g u r a t i o n e n . 
 
 V � l j   ' A n v � n d '   f � r   a t t   s t a r t a   o m   W i n S C P   m e d   e n   k o n f i g u r a t i o n   l a d d a d   f r � n   d e n   v a l d a   I N I - f i l e n .   D i n   n u v a r a n d e   k o n f i g u r a t i o n   k o m m e r   a t t   b e v a r a s   o c h   d u   k a n   � t e r g �   t i l l   d e n ,   o m   d e t   b e h � v s . | & S k r i v   � v e r | & A n v � n d =* * V i l l   d u   s k r i v a   � v e r   e n   s k r i v s k y d d a d   I N I - f i l   ' % s '   f � r   a t t   s p a r a   d i n   n u v a r a n d e   k o n f i g u r a t i o n ? * * D e n   h � r   f r � g a n   b l i r   i f r � g a s a t t   n � r   d u   h � l l e r   n e d   S h i f t - t a n g e n t e n   m e d a n   W i n S C P   s t � n g s   o c h   d i n   I N I - f i l   � r   s k r i v s k y d d a d .   N o r m a l t   s k r i v s   i n t e   I N I - f i l e r   � v e r   o c h   i n g a   � n d r i n g a r   i   k o n f i g u r a t i o n e n   g � r   f � r l o r a d e   n � r   W i n S C P   s t � n g s . K A v s l u t a   s e s s i o n e n   ' % s '   o c h   s t � n g   a p p l i k a t i o n e n   u t a n   a t t   s p a r a   e n   a r b e t s y t a ?                          W I N _ I N F O R M A T I O N    I n g a   s k i l l n a d e r   h i t t a d e s .  � p p n a r   s e s s i o n   ' % s ' 
 % s ' V � n t a r   p �   a t t   d o k u m e n t e t   s k a   s t � n g a s . . .  % s   ( � v e r f � r   m e d   % s )  % s   ( f � r   � v e r f � r i n g )  L o k a l :   % s 
 F j � r r :   % s  & T o u c h  & K � r     1 % d   f e l   u p p s t o d   v i d   s e n a s t e   o p e r a t i o n e n .   V i s a   d e m ?  F e l   % d   a v   % d : 
 % s  D u   h a r   d e n   s e n a s t e   v e r s i o n e n .  N y   v e r s i o n   % s   h a r   s l � p p t s .  P a r a m e t e r v � r d e :  ' % s '   k o m m a n d o p a r a m e t r a r                      U R L :   P r o t o k o l l e t   % s  A n s l u t e r . . .  F r � g a  F e l  P r o m p t 	 V � n t a r . . .  T a & r / G Z i p . . .  & A r k i v n a m n :  & U n T a r / G Z i p . . .  P a c k a   & u p p   t i l l   k a t a l o g :    & G r e p . . .  & S � k   e f t e r   m � n s t e r :  % d   L � s e r   k a t a l o g  B e r � k n a r . . .  
   
 % s  & U p p g r a d e r a   ; F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s '   v a l d e s   a u t o m a t i s k t . 4 � t e r g �   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s ' . + � t e r g �   t i l l   s t a n d a r d � v e r f � r i n g s i n s t � l l n i n g .  R e g e l   f � r   a u t o m a t i s k t   v a l : 
 % s    A d   H o c  P a u s a  & I n t e r n   e d i t o r �A p p l i k a t i o n   s t a r t a d   f � r   a t t   � p p n a   f i l   ' % s '   s t � n g d e s   f � r   t i d i g t .   O m   d e n   i n t e   s t � n g d e s   a v   d i g ,   d e   k a n   b e r o   p �   a t t   a p p l i k a t i o n e n   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   a p p l i k a t i o n e n   s k i c k a r   d �   d e n   n y a   f i l e n   t i l l   b e f i n t l i g   a p p l i k a t i o n   o c h   s t � n g s   o m e d e l b a r t .   W i n S C P   k a n   s t � d j a   s � d a n a   a p p l i k a t i o n e r   e n d a s t   s o m   e x t e r n   e d i t o r . 
   
 O m   d u   v i l l   a n v � n d a   a p p l i k a t i o n e n   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g a   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r .   = R e d i g e r a   ( e x t e r n ) | R e d i g e r a   v a l d a   f i l e r   m e d   e x t e r n   e d i t o r   ' % s ' � *   m a t c h a r   a l l a   a n t a l   t e c k e n . 
 ?   m a t c h a r   e x a k t   e t t   t e c k e n . 
 [ a b c ]   m a t c h a r   e t t   t e c k e n   f r � n   u p p s � t t n i n g e n . 
 [ a - z ]   m a t c h a r   e t t   t e c k e n   i   i n t e r v a l l e t . 
 E x e m p e l :   * . h t m l ;   p h o t o ? ? . p n g > M a s k   k a n   u t � k a s   m e d   s � k v � g s m a s k . 
 E x e m p e l :   * / p u b l i c _ h t m l / * . h t m l �M � n s t e r : 
 ! !   e x p a n d e r a r   t i l l   u t r o p s t e c k e n 
 !   e x p a n d e r a r   t i l l   f i l n a m n 
 ! &   e x p a n d e r a r   t i l l   l i s t a   m e d   v a l d a   f i l e r   ( c i t a t i o n s t e c k e n ,   m e l l a n s l a g s s e p a r e r a d ) 
 ! /   e x p a n d e r a r   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! S   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s - U R L 
 ! @   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s v � r d n a m n 
 ! U   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s a n v � n d a r n a m n 
 ! P   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s l � s e n o r d 
 ! #   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   p o r t n u m m e r 
 ! N   e x p a n d e r a r   t i l l   a k t u e l l t   s e s s i o n s n a m n 
 ! ? p r o m p t [ \ ] ? d e f a u l t !   e x p a n d e r a r   t i l l   a n v � n d a r v a l t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v t   \   u n d v i k e r   e s c a p e ) 
 ! ` c o m m a n d `   e x p a n d e r a r   t i l l   u t d a t a   a v   l o k a l t   k o m m a n d o 
   
 L o k a l t   k o m m a n d o m � n s t e r : 
 ! ^ !   e x p a n d e r a r   t i l l   f i l n a m n   f r � n   l o k a l   p a n e l 
   
 E x e m p e l : 
 g r e p   " ! ? M � n s t e r : ? ! "   ! & A A l l a   � v e r f � r i n g a r   i   b a k g r u n d e n   s l u t f � r d e s .   A n s l u t n i n g   a v s l u t a d e s .   L � s n i n g   a v   f j � r r k a t a l o g   a v b r � t s . ( S y n k r o n i s e r a d   b l � d d r i n g   s a t t e s   % s . | p � | a v ' V i s n i n g   a v   d o l d a   f i l e r   s a t t e s   % s . | p � | a v G A u t o m a t i s k   u p p d a t e r i n g   a v   f j � r r k a t a l o g   e f t e r   o p e r a t i o n   s a t t e s   % s . | p � | a v 1 � v e r f � r i n g   i   b a k g r u n d e n   k r � v e r   d i n   u p p m � r k s a m h e t .  � v e r f � r i n g s k � n   � r   t o m . Z ! Y   � r 
 ! M   m � n a d 
 ! D   d a g 
 ! T   t i d 
 ! P   p r o c e s s   i d 
 ! @   v � r d n a m n 
 ! S   s e s s i o n s n a m n 
 E x e m p e l : C : \ ! S ! T . l o g K P a s s i v t   l � g e   m � s t e   v a r a   a k t i v e r a d   n � r   F T P   a n s l u t n i n g   g e n o m   p r o x y   h a r   v a l t s . L U p p d a t e r i n g s k o n t r o l l   f � r   a p p l i k a t i o n e n   � r   t e m p o r � r t   a v s t � n g d .   F � r s � k   s e n a r e .  & G �   t i l l  V a d   � r   n y t t      O p e r a t i o n e n   s l u t f � r d e s  & P r i n t  & A s s o c i e r a d   a p p l i k a t i o n  P �  A v  A u t o S * * H u v u d l � s e n o r d e t   h a r   � n d r a t s . * * 
 
 D i n a   l a g r a d e   l � s e n o r d   � r   s � k r a d e   m e d   A E S - c h i f f e r .  H u v u d l � s e n o r d e t   h a r   � n d r a t s . S * * D u   h a r   t a g i t   b o r t   h u v u d l � s e n o r d e t . * * 
 
 D i n a   l a g r a d e   l � s e n o r d   � r   i n t e   s � k r a   l � n g r e .  H u v u d l � s e n o r d :      K o m m e r   a t t   k o n t r o l l e r a   i g e n :   % s  S e n a s t e   s e s s i o n e r Q M a s k e r   s k i l j s   � t   m e d   s e m i k o l o n   e l l e r   k o m m a .   
 P l a c e r a   u t e s l u t n a   m a s k e r   e f t e r   p i p e . , M a s k s l u t   m e d   s n e d s t r e c k   v � l j e r   u t   k a t a l o g e r .   � > s t o r l e k   m a t c h a r   f i l   s o m   � r   s t � r r e   � n   s t o r l e k 
 < s t o r l e k   m a t c h a r   f i l   m i n d r e   � n   s t o r l e k 
 > y y y y - m m - d d   m a t c h a r   f i l   s o m   � n d r a t s   e f t e r   d e t   d a t u m e t 
 < y y y y - m m - d d   m a t c h a r   f i l   s o m   � n d r a t s   f � r e   d e t   d a t u m e t 
 E x e m p e l :   * . z i p > 1 G ;   < 2 0 1 2 - 0 1 - 2 1  S e   h j � l p   f � r   f l e r   a l t e r n a t i v .  U T F - 8 � * * F � l j a n d e   a n v � n d a r s t a t i s t i k s d a t a   s k i c k a s   a n o n y m t   t i l l   W i n S C P . * * 
 
 U n d e r   t i d e n   k a n   a n n a n   s t a t i s t i k   s a m l a s   i n ,   k o m   g � r n a   t i l l b a k a   s e n a r e   f � r   a t t   k o n t r o l l e r a   e l l e r   k o n s u l t e r a   h j � l p e n . \ D e t   f i n n s   i n g e n   d a t a   i n s a m l a d   f � r   a n v � n d a r s t a t i s t i k   � n n u .   F � r s � k   i g e n   s e n a r e   e l l e r   s e   H j � l p .  � p p n a   w e b b p l a t s k a t a l o g   ' % s '  � p p n a r   a r b e t s y t a   ' % s '  S e n a s t e   a r b e t s y t o r  M i n   a r b e t s y t a - A r b e t s y t a   ' % s '   k o m m e r   a t t   s p a r a s   a u t o m a t i s k t .  A r b e t s y t a :   % s � * * � v e r f � r i n g s b e k r � f t e l s e   a v s t � n g d * * 
 
 D u   h a r   v a l t   a t t   i n t e   v i s a   d i a l o g r u t a n   f � r   � v e r f � r i n g s a l t e r n a t i v   n � s t a   g � n g .   K l i c k a   h � r   f � r   a t t   � n g r a .  F � r i n s t � l l n i n g a r 	 A v s l u t a d e u % s 
 
 D e t   u p p s t o d   n � g r a   f e l   v i d   k r y p t e r i n g e n   a v   l � s e n o r d   m e d   h j � l p   a v   e t t   n y t t   h u v u d l � s e n o r d   e l l e r   d e k r y p t e r a   l � s e n o r d . � W i n S C P   � r   e n   p o p u l � r   g r a t i s   S F T P -   o c h   F T P - k l i e n t   f � r   W i n d o w s ,   e n   k r a f t f u l l   f i l h a n t e r a r e   s o m   f � r b � t t r a r   p r o d u k t i v i t e t e n .   D e n   s t � d e r   � v e n   A m a z o n   S 3 ,   F T P S ,   S C P   o c h   W e b D A V - p r o t o k o l l .   P o w e r - a n v � n d a r e   k a n   a u t o m a t i s e r a   W i n S C P   m e d   . N E T   a s s e m b l y . 	 L a d d a r . . . * % s 
 
 K l i c k a   h � r   f � r   a t t   s e   v a d   s o m   � r   n y t t . # % d   s l �   u p p   l � n k a r   o c h   l � s e r   k a t a l o g  K a n   i n t e   v i s a  A n v � n d n i n g : 5 N a m n   p �   w e b b p l a t s   e l l e r   d i r e k t   s e s s i o n s s p e c i f i k a t i o n . ; � p p n a   s e s s i o n   i   e t t   n y t t   f � n s t e r ,   � v e n   o m   % A P P %   k � r s   r e d a n . % � p p n a r   f j � r r f i l   i   d e n   i n t e r n a   e d i t o r . ) S y n k r o n i s e r a s   i n n e h � l l e t   i   t v �   k a t a l o g e r . - S t a r t a r   f u n k t i o n e n   h � l l   f j � r r k a t a l o g   a k t u e l l . / S t a r t a r   o p e r a t i o n   u t a n   a t t   v i s a   a l t e r n a t i v r u t a . @ K o n s o l   ( t e x t )   l � g e .   S t a n d a r d l � g e ,   n � r   d e n   a n r o p a s   m e d   % A P P % . c o m . b K � r   b a t c h s k r i p t f i l .   O m   s k r i p t e t   i n t e   s l u t a r   m e d   ' e x i t ' - k o m m a n d o t ,   n o r m a l t   i n t e r a k t i v t   l � g e   f � l j e r .  K � r   l i s t a   m e d   s k r i p t k o m m a n d o n . + S k i c k a r   l i s t a   m e d   p a r a m e t r a r   t i l l   s k r i p t e t . # S � k v � g   t i l l   k o n f i g u r a t i o n s   I N I - f i l . D K o n f i g u r e r a r   i n s t � l l n i n g a r   m e d   h j � l p   a v   R A W - f o r m a t   s o m   i   e n   I N I - f i l . f U p p d a t e r i n g s i n s t � l l n i n g a r   a v   w e b b p l a t s e r   s o m   m a t c h a r   e n   m a s k   m e d   h j � l p   a v   r a w - f o r m a t   s o m   i   e n   I N I - f i l . # A k t i v e r a r   s e s s i o n l o g g n i n g   t i l l   f i l . E L o g g i n g s n i v �   ( 0 . . 2 ) ,   l � g g a   t i l l   *   f � r   a t t   a k t i v e r a   l � s e n o r d s l o g g n i n g .   A k t i v e r a r   X M L - l o g g n i n g   t i l l   f i l . 8 G r u p p e r a   a l l a   X M L - l o g e l e m e n t   s o m   t i l l h � r   s a m m a   k o m m a n d o .  S S H   p r i v a t   n y c k e l f i l ) F i n g e r a v t r y c k   a v   s e r v e r n s   S S H - v � r d n y c k e l .  T L S / S S L - k l i e n t c e r t i f i k a t f i l .  P a s s i v t   l � g e   ( F T P - p r o t o k o l l ) . ! I m p l i c i t   T L S / S S L   ( F T P - p r o t o k o l l ) . ! E x p l i c i t   T L S / S S L   ( F T P - p r o t o k o l l ) .  S e r v e r n   s v a r a d e   m e d   t i m e o u t . Q K o n f i g u r e r a r   a l l a   s e s s i o n s i n s t � l l n i n g a r   m e d   h j � l p   a v   R A W - f o r m a t   s o m   i   e n   I N I   f i l . + H e m s i d a   f � r   f � r f r � g n i n g a r   o m   u p p d a t e r i n g a r .  S k r i v e r   u t   d e n n a   a n v � n d n i n g . � K o n v e r t e r a r   p r i v a t   n y c k e l   t i l l   . p p k - f o r m a t   e l l e r   r e d i g e r a r   n y c k e l n .   A n v � n d   % s   f � r   a t t   a n g e   u t d a t a f i l .   A n v � n d   % s   f � r   a t t   � n d r a   e l l e r   s t � l l a   i n   l � s e n o r d s f r a s .   A n v � n d   % s   f � r   a t t   � n d r a   e l l e r   s t � l l a   i n   k o m m e n t a r e r . $ A n g e   l � s e n f r a s   f � r   a t t   s p a r a   n y c k e l : ) M a t a   � t e r   i n   l � s e n o r d s f r a s   f � r   v e r i f i e r a :  N y c k e l   s p a r a d   t i l l   " % s " . D F i n g e r a v t r y c k   f � r   s e r v e r   T L S / S S L - c e r t i f i k a t   ( e n d a s t   F T P S - p r o t o k o l l ) .  G e r   e t t   n a m n   t i l l   s e s s i o n e n � U p p d a t e r a r   f j � r r p a n e l e n   f � r   a l l a   i n s t a n s e r   a v   W i n S C P .   O m   e n   s e s s i o n   ( o c h   e v e n t u e l l t   e n   s � k v � g )   a n g e s ,   u p p d a t e r a r   e n d a s t   i n s t a n s e n   m e d   d e n   s e s s i o n e n   ( o c h   s � k v � g e n ) . ? A k t i v e r a r   l o g g r o t a t i o n   o c h   e v e n t u e l l t   r a d e r i n g   a v   g a m l a   l o g g a r .  L � s e n o r d e t   h a r   � n d r a t s .  � p p n a   & m � l m a p p e n  � p p n a   & n e d l a d d a d   f i l � * * K r y p t e r i n g s n y c k e l   g e n e r e r a d e s . * * 
 
 D u   b � r   s � k e r h e t s k o p i e r a   d e n   g e n e r e r a d e   k r y p t e r i n g s n y c k e l n .   O m   d u   f � r l o r a r   d e n   k a n   d u   i n t e   l � s a   d i n a   k r y p t e r a d e   f i l e r . > � p p n a   p l a t s p r o f i l   " % s " . | L o k a l   k a t a l o g : 
     % s | F j � r r k a t a l o g : 
     % s : S k r i v e r   u t   e n   l i s t a   � v e r   c h i f f e r   o c h   a l g o r i t m e r   s o m   s t � d s . H K o n f i g u r e r a r   � v e r f � r i n g s i n s t � l l n i n g a r   m e d   e t t   r � f o r m a t   s o m   i   e n   I N I - f i l . D ! E   e x p a n d e r a r   t i l l   s e r i a l i s e r a d e   a n s l u t n i n g s d a t a   f � r   a k t u e l l   s e s s i o n   F E t t   l � s e n o r d   f � r   e n   k r y p t e r a d   p r i v a t   n y c k e l   e l l e r   e t t   k l i e n t c e r t i f i k a t B T r y c k   p �   ' N e j '   f � r   a t t   a k t i v e r a   a u t o m a t i s k   s p a r n i n g   a v   a r b e t s y t a n . ( V � l j e r   d e n   a n g i v n a   f i l e n   i   f i l p a n e l e r n a . � * * R e d i g e r a   t e r m i n a l i n s t � l l n i n g a r   i   P u T T Y . * * 
 
 P u T T Y   k o m m e r   a t t   s t a r t a s .   R e d i g e r a   t e r m i n a l i n s t � l l n i n g a r   f � r   e n   t i l l f � l l i g   w e b b p l a t s   % s .   W i n S C P   k o m m e r   i h � g   d e s s a   i n s t � l l n i n g a r   e f t e r   a t t   d u   s t � n g e r   P u T T Y .  T e r m i n a l i n s t � l l n i n g a r   f � r   % s 8 E t t   a l t e r n a t i v t   s � t t   a t t   t i l l h a n d a h � l l a   e t t   a n v � n d a r n a m n 4 E t t   a l t e r n a t i v t   s � t t   a t t   t i l l h a n d a h � l l a   e t t   l � s e n o r d ! A l l a   p r o m p t e r   a v b r y t s   a u t o m a t i s k t R T i l l � t e r   s t r e a m i n g   a v   f i l e r   t i l l   s t d o u t   ( o c h   o m d i r i g e r a r   s t a t u s u t d a t a   t i l l   s t d e r r ) & T i l l � t e r   s t r � m n i n g   a v   f i l e r   f r � n   s t d i n                W I N _ F O R M S _ S T R I N G S          % s   f i l   ' % s '   t i l l   % s :  % s   % d   f i l e r   t i l l   % s :      l o k a l   k a t a l o g  f j � r r k a t a l o g    F l y t t a 	 s l � p p   m � l            T a r   b o r t  S t � l l e r   i n   i n s t � l l n i n g a r  T e m p o r � r   k a t a l o g 
 N y   k a t a l o g     	 A v m a r k e r a  M a r k e r a  % d   f i l  % d   f i l e r 
 % d   k a t a l o g  % d   k a t a l o g e r  % d   s y m b o l i s k   l � n k  % d   s y m b o l i s k a   l � n k a r    % s   E g e n s k a p e r  % s ,   . . .   E g e n s k a p e r  A n g e   g i l t i g t   g r u p p n a m n .  A n g e   g i l t i g t   � g a r n a m n .  T i l l b a k a   t i l l   % s  F r a m � t   t i l l   % s      A n s l u t n i n g s t i d  K o m p r i m e r i n g   ( % s )      I n f o r m a t i o n   o m   v a l d   f i l     P � p p n a   s p a r a d   s e s s i o n   ' % s '   ( h � l l   n e r e   S H I F T   f � r   a t t   � p p n a   s e s s i o n   i   n y t t   f � n s t e r )    L i c e n s   f � r   % s                � p p n a   k a t a l o g  H a n t e r a   b o k m � r k e n             
 R a d :   % d / % d 
 K o l u m n :   % d  T e c k e n :   % d   ( 0 x % . 2 x )  � n d r a d  K a n   i n t e   h i t t a   s t r � n g e n   ' % s ' .  T o t a l t   a n t a l   e r s � t t n i n g a r :   % d  G �   t i l l   r a d 
 R a d n u m m e r :  O g i l t i g t   r a d n u m m e r .  R e d i g e r a   l � n k / g e n v � g  L � g g   t i l l   l � n k / g e n v � g  I n t e   a n s l u t e n  A n s l u t e r . . .  V � l j   s e s s i o n   ' % s '  L � g g   t i l l   p l a t s p r o f i l  P l a t s p r o f i l n a m n :  F l y t t a   p l a t s p r o f i l  N y t t   k a t a l o g n a m n :  S p a r a   s e s s i o n   s o m  & S p a r a   s e s s i o n   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e )    K � r   e g e t   k o m m a n d o               5 % s ,   % d   p t 
 T h e   Q u i c k   B r o w n   F o x   J u m p s   O v e r   T h e   L a z y   D o g  O k � n d  B e r � k n a   k a t a l o g s t o r l e k        A l l m � n n a   i n s t � l l n i n g a r  L a g r a d e   s e s s i o n e r 
 C a c h e m i n n e  K o n f i g u r a t i o n e n s   I N I - f i l  S l u m p t a l s f r �   f i l  V � l j   l o k a l   k a t a l o g .  F l y t t a r      F l y t t a  H � l l   f j � r r k a t a l o g e n   u p p d a t e r a d % B e h � l l e r   f j � r r k a t a l o g e n   u p p d a t e r a d . . .  T e m p o r � r a   k a t a l o g e r  N y   f i l  R e d i g e r a   f i l  & S k r i v   f i l n a m n : ( D u p l i c a t e   f i l e   ' % s '   t o   r e m o t e   d i r e c t o r y : ' D u p l i c a t e   % d   f i l e s   t o   r e m o t e   d i r e c t o r y :  D u b b l e r a  K o p i e r a r  L � g g   t i l l   e g e t   k o m m a n d o  R e d i g e r a   e g e t   k o m m a n d o  L  F          H � & m t a   f l e r . . .  V � l j   e d i t o r a p p l i k a t i o n . 0 K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s   i   % s   a v   % s , L � g g   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g + R e d i g e r a   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g 	 S & t a n d a r d  & K o n f i g u r e r a . . .  E g & e t . . .  E g e t   k o m m a n d o  L � g g   t i l l   e d i t o r  R e d i g e r a   e d i t o r  % s ,   B a s e r a s   p �   % s   v e r s i o n   % s  & � p p n a    E n d a s t   & s a m m a   s t o r l e k   N u m b e r   o f   L i c e n s e s :   % s | U n l i m i t e d  P r o d u c t   I D :   % s  % s   ( E x p i r a t i o n   o n   % s )  % s       E d u c a t i o n a l   L i c e n s e  H � m t a r   e g e n s k a p e r    S S H   i m p l e m e n t a t i o n  K r y p t e r i n g s a l g o r i t m  K o m p r i m e r i n g  F i l � v e r f � r i n g s p r o t o k o l l  K a n   � n d r a   r � t t i g h e t e r  K a n   � n d r a   � g a r e / g r u p p  K a n   k � r a   g o d t y c k l i g t   k o m m a n d o " K a n   s k a p a   s y m b o l i s k   l � n k / h � r d   l � n k  K a n   s l �   u p p   a n v � n d a r g r u p p e r  K a n   d u b b l e r a   f j � r r f i l e r   $ � v e r f � r i n g s l � g e   f � r   r e n   t e x t   ( A S C I I ) $ K a n   k o n t r o l l e r a   t i l l g � n g l i g t   u t r y m m e  T o t a l t   a n t a l   b y t e s   p �   e n h e t  L e d i g t   a n t a l   b y t e s   p �   e n h e t   T o t a l t   a n t a l   b y t e s   f � r   a n v � n d a r e  L e d i g a   b y t e s   f � r   a n v � n d a r e  B y t e s   p e r   a l l o k e r i n g s e n h e t  O k � n d " H i t t a   P u T T Y / T e r m i n a l k l i e n t   k � r b a r a P P u T T Y / T e r m i n a l k l i e n t   k � r b a r a | % s | K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s | N / A  J � m f � r  S y n k r o n i s e r a r  A u t e n t i s e r i n g s b a n e r * I N I - f i l   ( * . i n i ) | * . i n i | A l l a   f i l e r   ( * . * ) | * . * ) V � l j   f i l   a t t   e x p o r t e r a   i n s t � l l n i n g a r   t i l l  S & e n a s t e :   % s  S & e n a s t e  B e r � k n a r   f i l k o n t r o l l s u m m a  K a n   b e r � k n a   f i l k o n t r o l l s u m m a  O k � n d  P r o t o k o l l   s o m   a n v � n d s    O s � k e r   a n s l u t n i n g  S � k e r   a n s l u t n i n g   ( % s )  E n d a s t   p r o t o k o l l k o m m a n d o n  F j � r r s y s t e m  K r y p t o g r a f i s k t   p r o t o k o l l      M i n a   d o k u m e n t 	 S k r i v b o r d    K o m m a n d o  S � t t   t i l l   s & t a n d a r d  - -   v a r n a   e f t e r   d e t t a   - -  3 D E S  B l o w f i s h  A E S  D E S  A r c f o u r  C h a C h a 2 0  - -   v a r n a   e f t e r   d e t t a   - -  D i f f i e - H e l l m a n   g r u p p   1  D i f f i e - H e l l m a n   g r u p p   1 4  D i f f i e - H e l l m a n   g r u p p   u t b y t e  R S A - b a s e r a t   n y c k e l u t b y t e  E C D H   n y c k e l u t b y t e  V � l j   l o k a l   p r o x y a p p l i k a t i o n � M � n s t e r : 
 \ n   f � r   n y   r a d 
 \ r   f � r   v a g n r e t u r 
 \ t   f � r   t a b b 
 \ x X X   f � r   h e x a d e c i m a l   a s c i i k o d 
 \ \   f � r   b a c k s l a s h 
 % v � r d   u t � k a s   t i l l   v � r d n a m n 
 % p o r t   u t � k a s   t i l l   p o r t n u m m e r 
 % u a n v � n d a r e   u t � k a s   t i l l   p r o x y a n v � n d a r n a m n 
 % l � s e n   u t � k a s   t i l l   p r o x y l � s e n o r d 
 % %   f � r   p r o c e n t t e c k e n = W e b b p l a t s k a t a l o g   e l l e r   a r b e t s y t a   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . E � r   d u   s � k e r   a t t   d u   v i l l   r a d e r a   s e s s i o n s k a t a l o g   ' % s '   m e d   % d   s e s s i o n e r ? $ K a n   i n t e   r a d e r a   s p e c i a l s e s s i o n   ' % s ' .  S k a p a   s e s s i o n s k a t a l o g  N y t t   k a t a l o g n a m n :    H o w   t o   p u r c h a s e   a   l i c e n s e . . .  M � l f j � r r & s � k v � g : � * * V i l l   d u   � p p n a   e n   s e p a r a t   s k a l s e s s i o n   f � r   a t t   d u b b l e r a   f i l e n ? * * 
 
 A k t u e l l   s e s s i o n   s t � d e r   i n t e   d i r e k t   d u b b l e r i n g   a v   f j � r r f i l e r .   S e p a r a t a   s k a l s e s s i o n e r   k a n   � p p n a s   f � r   a t t   b e a r b e t a   d u b b l e r i n g e n .   A l t e r n a t i v t   k a n   d u   d u b b l e r a   f i l e n   v i a   e n   l o k a l   t e m p o r � r   k o p i a .  E d i t o r    % s   d o l d  % s   f i l t r e r a d  F i l t e r � A k t u e l l   s e s s i o n   t i l l � t e r   e n d a s t   f � r � n d r i n g   a v   U I D   � g a n d e t .   D e t   v a r   i n t e   m � j l i g t   a t t   l � s a   U I D   f r � n   k o n t o n a m n e t   " % s " .   S p e c i f i c e r a   U I D   e x p l i c i t   i s t � l l e t .    � v e r f � r   i   & b a k g r u n d e n  % s   ( l � g g   t i l l   i   � v e r f � r i n g s k � )  I n g e n  V � l j   k o r t k o m m a n d o  K o r & t k o m m a n d o : 
 O b e g r � n s a t  H u v u d l � s e n o r d  & N u v a r a n d e   h u v u d l � s e n o r d :  N & y t t   h u v u d l � s e n o r d :  U p p r e p a   h u v u d l � s e n o r d : - S p a r a   & l � s e n o r d   ( s k y d d a s   g e n o m   h u v u d l � s e n o r d ) 	 L e t a   i   % s  S � k 	 S � k e r   . . .  K l a r . 	 A v b r u t e n .    & S t a r t  & S t o p p  S p a r a   & l � s e n o r d  A v b r y t e r . . .  K o d n i n g :   % s c F i l e n   h a r   � n d r a t s .   � n d r i n g a r   k o m m e r   a t t   g �   f � r l o r a d e ,   o m   f i l e n   l a d d a s   m e d   a n n a n   k o d n i n g .   F o r t s � t t a ? F � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   a r b e t s y t a n   ' % s '   m e d   % d   s e s s i o n ( e r ) ?    S p a r a   a r b e t s y t a   s o m  & S p a r a   a r b e t s y t a   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e ) . S p a r a   & l � s e n o r d   ( s o m   s k y d d a s   a v   h u v u d l � s e n o r d )  S p a r a   & l � s e n o r d Q � p p n a   a r b e t s y t a   ' % s '   ( h � l l   n e r   S h i f t   f � r   a t t   � p p n a   a r b e t s y t a n   i   e t t   n y t t   f � n s t e r )  & � p p n a   k a t a l o g U � p p n a   w e b b p l a t s k a t a l o g   ' % s '   ( h � l l   n e r   S h i f t   f � r   a t t   � p p n a   k a t a l o g   i   e t t   n y t t   f � n s t e r )    & S k a p a   g e n v � g   p �   s k r i v b o r d e t , A k t i v e r a   & a u t o m a t i s k t   s p a r a n d e   a v   a r b e t s y t a n  H � m t a  � v e r f � r  H � m t a  � v e r f � r ) % s   f i l   ' % s '   t i l l   % s   o c h   t a   b o r t   o r i g i n a l : + % s   % d   f i l e r   t i l l   % s   o c h   t a   b o r t   o r i g i n a l e n :  H � m t a   o c h   t a   b o r t  � v e r f � r   o c h   t a   b o r t  K �  I m p o r t e r a   w e b b p l a t s e r - F e l   v i d   l a d d n i n g   a v   f i l   ' % s '   m e d   ' % s '   k o d n i n g                        F e l   v i d   l a d d n i n g   a v   f i l   ' % s ' .  � t e r g � r   t i l l   ' % s '   k o d n i n g . ) V � l j   f i l   a t t   i m p o r t e r a   k o n f i g u r a t i o n   f r � n  S � k :   % s  ( t r y c k   p �   t a b b   f � r   n � s t a )  � v e r f � r  H � m t a r  % d   i   k � �M � n s t e r : 
 ! !   e x p a n d e r a r   t i l l   u t r o p s t e c k e n 
 ! /   e x p a n d e r a r   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! @   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   v � r d n a m n 
 ! U   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   a n v � n d a r n a m n 
 ! P   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   l � s e n o r d 
 ! #   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   p o r t n u m m e r 
 ! N   e x p a n d e r a r   t i l l   a k t u e l l t   s e s s i o n s n a m n 
 ! ? p r o m p t [ \ ] ? d e f a u l t !   e x p a n d e r a r   t i l l   a n v � n d a r v a l t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v t   \   u n d v i k e r   e s c a p e ) 
 ! ` c o m m a n d `   e x p a n d e r a r   t i l l   u t d a t a   a v   l o k a l t   k o m m a n d o  N y   w e b b p l a t s  K a t a l o g   w e b b p l a t s 	 A r b e t s y t a 8 D u   r e d i g e r a r   e n   w e b b p l a t s .   V i l l   d u   s p a r a   d i n a   � n d r i n g a r ? 	 & K a t a l o g :  < i n g e n >  S k a l  S C P / S k a l  E d i t o r  & I n g e n   f � r g 2 � t e r s t � l l   s e s s i o n   ( p a n e l )   f � r g   t i l l   s y s t e m s t a n d a r d  F & l e r   f � r g e r . . .  V � l j   f � r g   p �   s e s s i o n   ( p a n e l )  A & v l � g s n a   B O M   o c h   E O F   t e c k e n  A & v l � g s n a   B O M   t e c k e n   T L i c e n s a v t a l e n   f � r   f � l j a n d e   p r o g r a m   ( b i b l i o t e k )   � r   d e l   a v   a p p l i k a t i o n e n s   l i c e n s a v t a l .  V i s a   l i c e n s  T o o l b a r 2 0 0 0   l i b r a r y   % s  C o p y r i g h t   �   J o r d a n   R u s s e l l ! h t t p s : / / j r s o f t w a r e . o r g / t b 2 k d l . p h p  T B X   l i b r a r y   % s , C o p y r i g h t   �   A l e x   A .   D e n i s o v   a n d   c o n t r i b u t o r s ! h t t p s : / / g i t h u b . c o m / p l a s h e n k o v / T B X ' F i l e m a n a g e r   T o o l s e t   l i b r a r y   V e r s i o n   2 . 6  C o p y r i g h t   �   I n g o   E c k e l  J E D I   C o d e   L i b r a r y   ( J C L )   % s  h t t p s : / / j c l . d e l p h i - j e d i . o r g /  P n g C o m p o n e n t s   1 . 4 . 1 & C o p y r i g h t   �   U w e   R a a b e   a n d   M a r t i j n   S a l y ) h t t p s : / / g i t h u b . c o m / U w e R a a b e / P n g C o m p o n e n t s 	 S p a r a r . . .    S v e n s k   � v e r s � t t n i n g :  C o p y r i g h t   % s  F i l :  S � k v � g :  L � s n i n g 
 U p p l � s n i n g 	 & S t a n d a r d % � t e r s t � l l   e d i t o r n s   f � r g   t i l l   s t a n d a r d  V � l j   n � g o n   f � r g   t i l l   e d i t o r n  S p a r a   k o n v e r t e r a d   p r i v a t   n y c k e l ; P u T T Y   p r i v a t   n y c k e l f i l e r   ( * . p p k ) | * . p p k | A l l a   f i l e r   ( * . * ) | * . * / P r i v a t   n y c k e l   k o n v e r t e r a d   o c h   s p a r a d   t i l l   ' % s ' .    S k a p a   f i l - U R L  S k a p a   s e s s i o n - U R L / k o d  U R L  S k r i p t  k o d  D i t t   k o m m a n d o   % d  T i p s   % d   a v   % d  T i p s % K � r   a n p a s s a d e   k o m m a n d o t   ' % s '   s o m   ' % s '  K o m m a n d o r a d s a r g u m e n t  K o m m a n d o r a d s a r g u m e n t   f � r   % s K E n   s e r v e r v � r d s n y c k e l   � r   o k � n d .   A n s l u t   m i n s t   e n   g � n g ,   i n n a n   d u   s k a p a r   k o d e n .  C : \ s k r i v b a r \ s � k v � g \ t i l l \ l o g g \  S k a p a   & k o d . . .  S k a p a   � v e r f � r i n g s k o d   " K � r   s k r i p t e t   m e d   e t t   k o m m a n d o   s o m :   C : \ s � k v � g \ t i l l \ s c r i p t \ s c r i p t . t x t  D i n   k o d   ! K o n f i g u r e r a   � v e r f � r i n g s a l t e r n a t i v  � v e r f � r   f i l e r c E t t   t e s t f i l l i s t a   a n v � n d s   e n d a s t ,   � v e r v � g   a t t   a n v � n d a   e n   f i l m a s k   f � r   a t t   v � l j a   f i l e r   f � r   � v e r f � r i n g .  S � k   e f t e r   u p p d a t e r i n g a r  L � g g   t i l l   u t � k n i n g $ A n g e   U R L   e l l e r   s � k v � g   t i l l   u t � k n i n g :     
 B l � d d r a . . . 	 V � l j   ' % s '  & P a u s a   i   s l u t e t  & S e s s i o n s l o g g f i l  V � l j   f i l   f � r   s e s s i o n s l o g g . 4 S e s s i o n s l o g g f i l a r   ( * . l o g ) | * . l o g | A l l a   f i l e r   ( * . * ) | * . *  A n v � n d a r s t a t i s t i k    & F i l t e r :  & K o p i e r a   t i l l   u r k l i p p  V � r d :   % s 
 V � r d n y c k e l :   % s  K & o p i e r a  & M a r k e r a   a l l t  K o r & t k o m m a n d o :                    A l l m � n t  A n s l u t e n 0 A n s l u t e n   m e d   % s .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .   * A n s l u t e n   m e d   % s ,   f � r m e d l a r   S S L - k o p p l i n g . . .  A n s l u t e r   t i l l   % s   . . .  L i s t n i n g   a v   k a t a l o g e r   l y c k a d  K o p p l a r   i f r � n   s e r v e r    s t a r t a r   n e r l a d d n i n g   a v   % s  N e r l a d d n i n g   l y c k a d   * F � r s � k e r   a t t   a n s l u t a   % s   g e n o m   F T P   p r o x y . . .                 � t e r f � r   l i s t n i n g   a v   k a t a l o g e r . . . 7 S S L - k o p p l i n g   u p p r � t t a d .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .  S S L - k o p p l i n g   u p p r � t t a d  S t a r t a r   � v e r f � r i n g   a v   % s  � v e r f � r i n g   l y c k a d     # H � m t a r   f i l i n f o r m a t i o n   f r a m g � n g s r i k t  H � m t a r   f i l i n f o r m a t i o n . . .  K u n d e   i n t e   h � m t a   f i l i n f o r m a t i o n                   5 K u n d e   i n t e   s k a p a   s o c k e t   i   d e n   a n g i v n a   p o r t i n t e r v a l l e t    K a n   i n t e   u p p r � t t a   S S L - k o p p l i n g   ' K u n d e   i n t e   � t e r f �   l i s t n i n g   a v   k a t a l o g e r     # K a n   i n t e   i n i t i a l i s e r a   S S L - b i b l i o t e k         , � v e r f � r i n g s t u n n e l   k a n   i n t e   � p p n a s .   O r s a k :   % s    K a n   i n t e   t o l k a   v � r d n a m n   " % s " > � t e r u p p t a g n i n g s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   s k r i v a   � v e r   f i l . I P a u s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   m e n   l o k a l   o c h   f j � r r f i l s t o r l e k   � r   l i k a . , O f � r m � g e n   a t t   s k i c k a   k o m m a n d o .   K o p p l a   i f r � n .    P e e r   c e r t i f i k a t   f � r k a s t a s    N e r l a d d n i n g   a v b r u t e n                      F i l e n   f i n n s   r e d a n          P r o x y   k r � v e r   a u t e n t i s e r i n g P N � d v � n d i g   a u t e n t i s e r i n g s t y p   r a p p o r t e r a d   a v   p r o x y s e r v e r   � r   o k � n d   e l l e r   s t � d s   i n t e % K a n   i n t e   a v g � r a   v � r d   t i l l   p r o x y s e r v e r ! K a n   i n t e   a n s l u t a   t i l l   p r o x y s e r v e r C B e g � r a n   f r � n   p r o x y   m i s s l y c k a d e s ,   k a n   i n t e   a n s l u t a   g e n o m   p r o x y s e r v e r                        T i m e o u t   d e t e k t e r a d .  � v e r f � r i n g   a v b r u t e n            K u n d e   i n t e   s � t t a   f i l p e k a r e  O k � n t   f e l   i   S S L - l a g r e t % K u n d e   i n t e   v e r i f i e r a   S S L - c e r t i f i k a t e t                                                            1 0 0     5 A n s l u t n i n g   m e d   p r o x y   e t a b l e r a d ,   u t f � r   h a n d s k a k n i n g . . .  k o n t r o l l a n s l u t n i n g  d a t a a n s l u t n i n g                            W I N _ V A R I A B L E $ C o p y r i g h t   �   2 0 0 0  2 0 2 2   M a r t i n   P r i k r y l  h t t p s : / / w i n s c p . n e t / # h t t p s : / / w i n s c p . n e t / e n g / d o c s / h i s t o r y    h t t p s : / / w i n s c p . n e t / f o r u m /  h t t p s : / / w i n s c p . n e t / u p d a t e s . p h p # h t t p s : / / w i n s c p . n e t / e n g / d o w n l o a d . p h p ! h t t p s : / / w i n s c p . n e t / e n g / d o n a t e . p h p + h t t p s : / / w i n s c p . n e t / e n g / d o c s / ? v e r = % s & l a n g = % s - h t t p s : / / w i n s c p . n e t / e n g / d o c s / % s ? v e r = % s & l a n g = % s ' h t t p s : / / w i n s c p . n e t / e n g / t r a n s l a t i o n s . p h p : h t t p s : / / w i n s c p . n e t / e n g / d o c s / s e a r c h . p h p ? v e r = % s & l a n g = % s & q = % s K h t t p s : / / w i n s c p . n e t / f o r u m / p o s t i n g . p h p ? m o d e = n e w t o p i c & v e r = % s & l a n g = % s & r e p o r t = % s " h t t p s : / / w i n s c p . n e t / e n g / u p g r a d e . p h p 8 h t t p s : / / w w w . m i c r o s o f t . c o m / s t o r e / a p p s / 9 p 0 p q 8 b 6 5 n 8 x ? c i d = % s   + h t t p s : / / w i n s c p . n e t / e n g / d o c s / m i c r o s o f t _ s t o r e 1 h t t p s : / / w i n s c p . n e t / u p d a t e n e w s . p h p ? s t o r e _ g e t _ i m g = 1                                             5 G e n e r a t e H t t p U r l . G e n e r a t e   & H T T P   U R L = G e n e r e r a   & H T T P - U R L ^ G e n e r a t e H t t p U r l . G e n e r a t e s   H T T P   U R L   o f   t h e   s e l e c t e d   f i l e = G e n e r e r a r   H T T P - U R L   f � r   d e n   v a l d a   f i l e n  G e n e r a t e H t t p U r l . U R L = U R L T G e n e r a t e H t t p U r l . T h e s e   o p t i o n s   a r e   s i t e - s p e c i f i c . = D e s s a   a l t e r n a t i v   � r   p l a t s s p e c i f i k a . 8 G e n e r a t e H t t p U r l . & W e b   r o o t   p a t h : = & W e b b s e r v e r n s   r o t s � k v � g : ( G e n e r a t e H t t p U r l . U s e   H T T P & S = A n v � n d   H T T P & S C G e n e r a t e H t t p U r l . & U R L   r o o t   p a t h   ( o p t i o n a l ) : = & U R L   r o t s � k v � g   ( v a l f r i ) : c G e n e r a t e H t t p U r l . & W e b   s e r v e r   h o s t n a m e   o v e r r i d e   ( o p t i o n a l ) : = � s i d o s � t t   w e b b s e r v e r n s   v � r d n a m n   ( v a l f r i ) : " G e n e r a t e H t t p U r l . O p t i o n s = A l t e r n a t i v $ G e n e r a t e H t t p U r l . D i s p l a y   U R L = V i s a   U R L > G e n e r a t e H t t p U r l . C o p y   U R L   t o   c l i p b o a r d = K o p i e r a   U R L   t i l l   u r k l i p p ? G e n e r a t e H t t p U r l . O p e n   U R L   i n   w e b   b r o w s e r = � p p n a   U R L   i   w e b b l � s a r e n ) C o m p a r e F i l e s . & C o m p a r e   F i l e s = & J � m f � r   f i l e r � C o m p a r e F i l e s . C o m p a r e s   t h e   s e l e c t e d   l o c a l   a n d   r e m o t e   p a t h   u s i n g   a n   e x t e r n a l   f i l e   c o m p a r i s o n   t o o l = J � m f � r   v a l d   l o k a l   o c h   f j � r r s � k v � g   m e d   h j � l p   a v   e t t   e x t e r n t   v e r k t y g   f � r   j � m f � r e l s e   a v   f i l e r  C o m p a r e F i l e s . O p t i o n s = A l t e r n a t i v C C o m p a r e F i l e s . S e l e c t   & f i l e   c o m p a r i s o n   t o o l : = V � l j   & j � m f � r e l s e v e r k t y g : ! C o m p a r e F i l e s . A u t o m a t i c = A u t o m a t i s k < V e r i f y F i l e C h e c k s u m . V e r i f y   & C h e c k s u m = V e r i f i e r a   & k o n t r o l l s u m m a � V e r i f y F i l e C h e c k s u m . C o m p a r e s   c h e c k s u m s   o f   t h e   s e l e c t e d   l o c a l   a n d   r e m o t e   f i l e = J � m f � r   k o n t r o l l s u m m o r   f � r   d e n   v a l d a   l o k a l a   o c h   f j � r r f i l e n 1 S e a r c h T e x t . & S e a r c h   f o r   T e x t . . . = & S � k   e f t e r   t e x t . . . � S e a r c h T e x t . S e a r c h e s   r e c u r s i v e l y   f o r   a   t e x t   i n   t h e   c u r r e n t   r e m o t e   d i r e c t o r y = S � k e r   r e k u r s i v t   e f t e r   e n   t e x t   i   d e n   a k t u e l l a   f j � r r k a t a l o g e n  S e a r c h T e x t . T e x t : = T e x t :  S e a r c h T e x t . F i l e   m a s k : = F i l m a s k : 2 Z i p U p l o a d . & Z I P   a n d   U p l o a d . . . = & Z I P   o c h   l a d d a   u p p . . .   � Z i p U p l o a d . P a c k s   t h e   s e l e c t e d   f i l e s   t o   a   Z I P   a r c h i v e   a n d   u p l o a d s   i t = P a k e t e r a r   d e   v a l d a   f i l e r n a   t i l l   e t t   Z I P - a r k i v   o c h   l a d d a r   u p p   d e t   $ Z i p U p l o a d . & A r c h i v e   n a m e : = & A r k i v n a m n : " Z i p U p l o a d . U s e   & 7 - z i p = A n v � n d   & 7 - z i p < Z i p U p l o a d . A r c h i v e   & t y p e   ( w i t h   7 - z i p ) : = A r k i v & t y p   ( m e d   7 - z i p ) : F Z i p U p l o a d . 7 - z i p   & p a t h   ( 7 z . e x e / 7 z a . e x e ) : = 7 - z i p   s � k v � g   ( 7 z . e x e / 7 z a . e x e ) :  Z i p U p l o a d . L o g g i n g = L o g g n i n g W K e e p L o c a l U p T o D a t e . & K e e p   L o c a l   D i r e c t o r y   u p   t o   D a t e . . . = & H � l l   l o k a l   k a t a l o g   u p p d a t e r a d . . . � K e e p L o c a l U p T o D a t e . P e r i o d i c a l l y   s c a n s   f o r   c h a n g e s   i n   a   r e m o t e   d i r e c t o r y   a n d   r e f l e c t s   t h e m   o n   a   l o c a l   d i r e c t o r y = S k a n n a r   p e r i o d i s k t   e f t e r   f � r � n d r i n g a r   i   e n   f j � r r k a t a l o g   o c h   � t e r s p e g l a r   d e m   p �   e n   l o k a l   k a t a l o g ' K e e p L o c a l U p T o D a t e . D i r e c t o r i e s = K a t a l o g e r h K e e p L o c a l U p T o D a t e . & W a t c h   f o r   c h a n g e s   i n   t h e   r e m o t e   d i r e c t o r y : = & T i t t a   e f t e r   f � r � n d r i n g a r   i   f j � r r k a t a l o g e n � K e e p L o c a l U p T o D a t e . . . .   & a n d   a u t o m a t i c a l l y   r e f l e c t   t h e m   o n   t h e   l o c a l   d i r e c t o r y : = . . .   & o c h   r e f l e k t e r a   d e m   a u t o m a t i s k t   p �   d e n   l o k a l a   k a t a l o g e n : $ K e e p L o c a l U p T o D a t e . O p t i o n s = A l t e r n a t i v . K e e p L o c a l U p T o D a t e . & D e l e t e   f i l e s = & T a   b o r t   f i l e r < K e e p L o c a l U p T o D a t e . & B e e p   o n   c h a n g e = & S y s t e m l j u d   v i d   f � r � n d r i n g 6 K e e p L o c a l U p T o D a t e . C o n t i n u e   o n   & e r r o r = F o r t s � t t   v i d   & f e l A K e e p L o c a l U p T o D a t e . & I n t e r v a l   ( i n   s e c o n d s ) : = I n t e r v a l l   ( i   s e k u n d e r ) : " K e e p L o c a l U p T o D a t e . L o g g i n g = L o g g n i n g 0 B a t c h R e n a m e . B a t c h   & R e n a m e . . . = B a t c h ,   & b y t   n a m n . . . w B a t c h R e n a m e . R e n a m e s   r e m o t e   f i l e s   u s i n g   a   r e g u l a r   e x p r e s s i o n = B y t e r   n a m n   p �   f j � r r f i l e r   m e d   h j � l p   a v   e t t   r e g u l j � r t   u t t r y c k  B a t c h R e n a m e . R e n a m e = B y t   n a m n j B a t c h R e n a m e . R e p l a c e   f i l e   n a m e   p a r t   m a t c h i n g   t h i s   p a t t e r n : = E r s � t t   d e l   a v   f i l n a m n   s o m   m a t c h a r   d e t t a   m � n s t e r :  B a t c h R e n a m e . w i t h : = m e d :  B a t c h R e n a m e . O p t i o n s = A l t e r n a t i v 4 B a t c h R e n a m e . & P r e v i e w   c h a n g e s = F � & r h a n d s v i s a   � n d r i n g a r  B a t c h R e n a m e . L o g g i n g = L o g g n i n g ? A r c h i v e D o w n l o a d . & A r c h i v e   a n d   D o w n l o a d . . . = & A r k i v e r a   o c h   h � m t a . . . A r c h i v e D o w n l o a d . P a c k s   t h e   s e l e c t e d   f i l e s   t o   a n   a r c h i v e ,   d o w n l o a d s   i t ,   a n d   o p t i o n a l l y   e x t r a c t s   t h e   a r c h i v e   t o   t h e   c u r r e n t   l o c a l   d i r e c t o r y = P a c k a r   d e   v a l d a   f i l e r n a   t i l l   e t t   a r k i v ,   l a d d a r   n e r   d e t   o c h   e x t r a h e r a r   e v e n t u e l l t   a r k i v e t   t i l l   d e n   a k t u e l l a   l o k a l a   k a t a l o g e n * A r c h i v e D o w n l o a d . & A r c h i v e   n a m e : = & A r k i v n a m n : ) A r c h i v e D o w n l o a d . A r c h i v e   & t y p e : = A r k i v & t y p :   A r c h i v e D o w n l o a d . P a c k i n g = P a c k n i n g A A r c h i v e D o w n l o a d . C u s t o m   a r c h i v e   & c o m m a n d : = A n p a s s a t   a r k i v & k o m m a n d o : % A r c h i v e D o w n l o a d . E x t r a c t i n g = U p p a c k n i n g @ A r c h i v e D o w n l o a d . & E x t r a c t   a f t e r   d o w n l o a d = & P a c k   u p p   e f t e r   h � m t n i n g F A r c h i v e D o w n l o a d . U s e   & 7 - z i p   f o r   e x t r a c t i n g = A n v � n d   & 7 - z i p   f � r   u p p a c k n i n g L A r c h i v e D o w n l o a d . 7 - z i p   & p a t h   ( 7 z . e x e / 7 z a . e x e ) : = 7 - z i p   s � k v � g   ( 7 z . e x e / 7 z a . e x e ) :   A r c h i v e D o w n l o a d . L o g g i n g = L o g g n i n g m S y n c h r o n i z e A n o t h e r S e r v e r . & S y n c h r o n i z e   w i t h   A n o t h e r   R e m o t e   S e r v e r . . . = & S y n k r o n i s e r a   m e d   e n   a n n a n   f j � r r s e r v e r . . . S y n c h r o n i z e A n o t h e r S e r v e r . S y n c h r o n i z e s   a   d i r e c t o r y   o n   a n o t h e r   s e r v e r   ( o r   a n o t h e r   d i r e c t o r y   o n   t h i s   s e r v e r )   a g a i n s t   a   d i r e c t o r y   o n   t h i s   s e r v e r = S y n k r o n i s e r a r   e n   k a t a l o g   p �   e n   a n n a n   s e r v e r   ( e l l e r   e n   a n n a n   k a t a l o g   p �   d e n   h � r   s e r v e r n )   m o t   e n   k a t a l o g   p �   d e n   h � r   s e r v e r n j S y n c h r o n i z e A n o t h e r S e r v e r . S y n c h r o n i z e   d i r e c t o r y   f r o m   & t h i s   s e r v e r : = S y n k r o n i s e r a   k a t a l o g   f r � n   & d e n n a   s e r v e r : . S y n c h r o n i z e A n o t h e r S e r v e r . & D i r e c t o r y : = & K a t a l o g : K S y n c h r o n i z e A n o t h e r S e r v e r . . . .   t o   & a n o t h e r   s e r v e r : = . . .   t i l l   e n   & a n n a n   s e r v e r : , S y n c h r o n i z e A n o t h e r S e r v e r . & S e s s i o n : = & S e s s i o n : Y S y n c h r o n i z e A n o t h e r S e r v e r . & P r o m p t   f o r   s e s s i o n   p a s s w o r d = & F r � g a   e f t e r   l � s e n o r d   f � r   s e s s i o n e n . S y n c h r o n i z e A n o t h e r S e r v e r . D i & r e c t o r y : = K a & t a l o g : + S y n c h r o n i z e A n o t h e r S e r v e r . O p t i o n s = A l t e r n a t i v 5 S y n c h r o n i z e A n o t h e r S e r v e r . & D e l e t e   f i l e s = & T a   b o r t   f i l e r A S y n c h r o n i z e A n o t h e r S e r v e r . & P r e v i e w   c h a n g e s = F � & r h a n d s v i s a   � n d r i n g a r = S y n c h r o n i z e A n o t h e r S e r v e r . C o n t i n u e   o n   & e r r o r = F o r t s � t t   v i d   & f e l   ) S y n c h r o n i z e A n o t h e r S e r v e r . L o g g i n g = L o g g n i n g                                 " S k a l t i l l � g g e t   � r   i n t e   i n s t a l l e r a t . 7 S k a l t i l l � g g e t   � r   i n s t a l l e r a t ,   m e n   d e t   h a r   i n t e   l a d d a t s . % S k a l t i l l � g g e t   i n s t a l l e r a s   o c h   l a d d a s . E * * P u b l i k   n y c k e l   f � r   a t t   k l i s t r a   i n   i   O p e n S S H   a u t h o r i z e d _ k e y s - f i l e n : * * � * * I n s t a l l e r a   d e n   p u b l i k a   n y c k e l n   t i l l   i c k e - O p e n S S H   s e r v e r ? * * 
 
 I n s t a l l e r i n g   a v   d e n   p u l i k a   n y c k e l n   s t � d s   e n d a s t   f � r   O p e n S S H   s e r v e r   ( a u t h o r i z e d _ k e y s - f i l ) . 
 
 D i n   s e r v e r   � r   % s . ! I n s t a l l e r a r   p u b l i k   n y c k e l   " % s " . . . U * * P u b l i k   n y c k e l   " % s "   i n s t a l l e r a d e s . * * 
 
 D u   k a n   n u   l o g g a   i n   p �   s e r v e r n   m e d   n y c k e l p a r e t . l E v e n t u e l l a   f e l   b e h � r i g h e t e r   f � r   f i l e n   " % s "   o c h / e l l e r   d e s s   f � r � l d r a m a p p   u p p t � c k t e s .   V � n l i g e n   k o n t r o l l e r a   d e m . * V � l j   n y c k e l   f � r   a t t   i n s t a l l e r a   t i l l   s e r v e r � P u T T Y   p r i v a t a   n y c k e l f i l e r   ( * . p p k ) | * . p p k | A l l a   p r i v a t a   n y c k e l f i l e r   ( * . p p k ; * . p e m ; * . k e y ; i d _ * ) | * . p p k ; * . p e m ; * . k e y ; i d _ * | A l l a   f i l e r   ( * . * ) | * . *  C h e c k l i s t   f � r   s y n k r o n i s e r i n g  S k r i v s k y d d a d  B e r � k n a r  S p a r a   s o m   & f � r i n s t � l l n i n g . . .  B y t   n a m n   p �   s e s s i o n  & N y t t   s e s s i o n s n a m n :  S y n k r o n i s e r i n g e n   s l u t f � r d e s . � U p p l a d d a d e   f i l e r :   % s   ( % s ) | N e d l a d d a d e   f i l e r :   % s   ( % s ) | L o k a l a   f i l e r   r a d e r a d e :   % s | E x t e r n a   f i l e r   r a d e r a d e :   % s | J � m f � r e l s e t i d :   % s | S y n k r o n i s e r i n g s t i d :   % s 1 S k a l t i l l � g g   k a n   i n t e   f u n g e r a   p �   d e t   h � r   s y s t e m e t .  F i l f � r g � F � r   a t t   a k t i v e r a   a u t o m a t i s k a   u p p d a t e r i n g a r ,   s n � l l a   < a   h r e f = " % D O N A T E _ U R L % " > d o n e r a   t i l l   W i n S C P - u t v e c k l i n g < / a >   e l l e r   % G E T _ I M G %   W i n S C P   f r � n   < a   h r e f = " % S T O R E _ U R L % " > M i c r o s o f t   S t o r e < / a > .  N y 	 S t a t i s t i k  R a w - w e b b p l a t s i n s t � l l n i n g a r  & L � g g   t i l l . . . " L � g g   t i l l   R a w - w e b b p l a t s i n s t � l l n i n g  & W e b b p l a t s i n s t � l l n i n g :  L a d d a   u p p   n y   l o k a l   f i l  L a d d a   n e r   n y   f j � r r f i l  L a d d a   u p p   u p p d a t e r a d   l o k a l   f i l  L a d d a   n e r   u p p d a t e r a d   f j � r r f i l  T a   b o r t   f � r � l d r a d   f j � r r f i l    T a   b o r t   f � r � l d r a d   l o k a l   f i l  K l i c k a   f � r   o m v � n t                                          a n   u n n a m e d   f i l e                      N o   e r r o r   m e s s a g e   i s   a v a i l a b l e . ' A n   u n s u p p o r t e d   o p e r a t i o n   w a s   a t t e m p t e d . $ A   r e q u i r e d   r e s o u r c e   w a s   u n a v a i l a b l e .  O u t   o f   m e m o r y .  A n   u n k n o w n   e r r o r   h a s   o c c u r r e d .                                        F a i l e d   t o   l a u n c h   h e l p .  I n t e r n a l   a p p l i c a t i o n   e r r o r .  C o m m a n d   f a i l e d . ) I n s u f f i c i e n t   m e m o r y   t o   p e r f o r m   o p e r a t i o n . P S y s t e m   r e g i s t r y   e n t r i e s   h a v e   b e e n   r e m o v e d   a n d   t h e   I N I   f i l e   ( i f   a n y )   w a s   d e l e t e d . B N o t   a l l   o f   t h e   s y s t e m   r e g i s t r y   e n t r i e s   ( o r   I N I   f i l e )   w e r e   r e m o v e d . F T h i s   p r o g r a m   r e q u i r e s   t h e   f i l e   % s ,   w h i c h   w a s   n o t   f o u n d   o n   t h i s   s y s t e m . t T h i s   p r o g r a m   i s   l i n k e d   t o   t h e   m i s s i n g   e x p o r t   % s   i n   t h e   f i l e   % s .   T h i s   m a c h i n e   m a y   h a v e   a n   i n c o m p a t i b l e   v e r s i o n   o f   % s .      P l e a s e   e n t e r   a n   i n t e g e r .  P l e a s e   e n t e r   a   n u m b e r . * P l e a s e   e n t e r   a n   i n t e g e r   b e t w e e n   % 1   a n d   % 2 . ( P l e a s e   e n t e r   a   n u m b e r   b e t w e e n   % 1   a n d   % 2 . ( P l e a s e   e n t e r   n o   m o r e   t h a n   % 1   c h a r a c t e r s .  P l e a s e   s e l e c t   a   b u t t o n . * P l e a s e   e n t e r   a n   i n t e g e r   b e t w e e n   0   a n d   2 5 5 .   P l e a s e   e n t e r   a   p o s i t i v e   i n t e g e r .   P l e a s e   e n t e r   a   d a t e   a n d / o r   t i m e .  P l e a s e   e n t e r   a   c u r r e n c y .                U n e x p e c t e d   f i l e   f o r m a t . V % 1 
 C a n n o t   f i n d   t h i s   f i l e . 
 P l e a s e   v e r i f y   t h a t   t h e   c o r r e c t   p a t h   a n d   f i l e   n a m e   a r e   g i v e n .  D e s t i n a t i o n   d i s k   d r i v e   i s   f u l l . 5 U n a b l e   t o   r e a d   f r o m   % 1 ,   i t   i s   o p e n e d   b y   s o m e o n e   e l s e . A U n a b l e   t o   w r i t e   t o   % 1 ,   i t   i s   r e a d - o n l y   o r   o p e n e d   b y   s o m e o n e   e l s e . . A n   u n e x p e c t e d   e r r o r   o c c u r r e d   w h i l e   r e a d i n g   % 1 . . A n   u n e x p e c t e d   e r r o r   o c c u r r e d   w h i l e   w r i t i n g   % 1 .                                           # U n a b l e   t o   r e a d   w r i t e - o n l y   p r o p e r t y . # U n a b l e   t o   w r i t e   r e a d - o n l y   p r o p e r t y .      N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  % 1   w a s   n o t   f o u n d .  % 1   c o n t a i n s   a n   i n v a l i d   p a t h . = % 1   c o u l d   n o t   b e   o p e n e d   b e c a u s e   t h e r e   a r e   t o o   m a n y   o p e n   f i l e s .  A c c e s s   t o   % 1   w a s   d e n i e d . . A n   i n v a l i d   f i l e   h a n d l e   w a s   a s s o c i a t e d   w i t h   % 1 . < % 1   c o u l d   n o t   b e   r e m o v e d   b e c a u s e   i t   i s   t h e   c u r r e n t   d i r e c t o r y . 6 % 1   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   t h e   d i r e c t o r y   i s   f u l l .  S e e k   f a i l e d   o n   % 1 5 A   h a r d w a r e   I / O   e r r o r   w a s   r e p o r t e d   w h i l e   a c c e s s i n g   % 1 . 0 A   s h a r i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . 0 A   l o c k i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  D i s k   f u l l   w h i l e   a c c e s s i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d .    N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . / A n   a t t e m p t   w a s   m a d e   t o   w r i t e   t o   t h e   r e a d i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d . 0 A n   a t t e m p t   w a s   m a d e   t o   r e a d   f r o m   t h e   w r i t i n g   % 1 .  % 1   h a s   a   b a d   f o r m a t . " % 1   c o n t a i n e d   a n   u n e x p e c t e d   o b j e c t .   % 1   c o n t a i n s   a n   i n c o r r e c t   s c h e m a .                 0 C a n n o t   c o n v e r t   s c i e n t i f i c   n o t a t i o n   t o   T B c d   v a l u e   C a n n o t   c o n v e r t   N A N   t o   T B c d   v a l u e ( I n v a l i d   B c d   P r e c i s i o n   ( % d )   o r   S c a l e   ( % d ) : C a n n o t   c o n v e r t   t o   T B c d :   s t r i n g   h a s   m o r e   t h a n   6 4   d i g i t s :   % s  % s   i s   n o t   a   v a l i d   h e x   s t r i n g  U n s u p p p o r t e d   v a r i a n t   t y p e   % d  v a r D i s p a t c h   t y p e   n o t   s u p p o r t e d  v a r E r r o r   t y p e   n o t   s u p p o r t e d  B C D   o v e r f l o w  % s   i s   n o t   a   v a l i d   B C D   v a l u e 2 I n v a l i d   H T M L   e n c o d e d   c h a r a c t e r   ( % s )   a t   p o s i t i o n   % d           & A t t e m p t i n g   t o   h o o k   c h i l d   w i n d o w s   t w i c e  S a v e   t h e   c u r r e n t   f i l e ? F I n t e r n a l   e r r o r :   d a t a   t y p e   k i n d   % s   c a n n o t   b e   c o n v e r t e d   t o   a n d   f r o m   t e x t + I n v o k a b l e   C l a s s   % s   i m p l e m e n t s   n o   i n t e r f a c e s  T y p e   c a n n o t   b e   c a s t   a s   V a r i a n t  I n t e r f a c e   % s   h a s   n o   R T T I 5 P a r a m e t e r   % s   o n   M e t h o d   % s   o f   I n t e r f a c e   % s   h a s   n o   R T T I  I n v a l i d   d a t e   s t r i n g :   % s  I n v a l i d   t i m e   s t r i n g :   % s  I n v a l i d   m i n u t e :   % d  I n v a l i d   m i l l i s e c o n d :   % d  I n v a l i d   f r a c t i o n a l   s e c o n d :   % f  I n v a l i d   h o u r   o f f s e t :   % d  I n v a l i d   d u r a t i o n   s t r i n g :   % s # H o u r   O f f s e t   p o r t i o n   o f   t i m e   i n v a l i d  I n v a l i d   d e c i m a l   s t r i n g :   ' ' % s ' '   D 3 r d - l e v e l   c a c h e :   1 8   M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 3 r d - l e v e l   c a c h e :   2 4   M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e  6 4 - B y t e   P r e f e t c h i n g  1 2 8 - B y t e   P r e f e t c h i n g e C P U I D   l e a f   2   d o e s   n o t   r e p o r t   c a c h e   d e s c r i p t o r   i n f o r m a t i o n ,   u s e   C P U I D   l e a f   4   t o   q u e r y   c a c h e   p a r a m e t e r s 	 W i n d o w s   8  W i n d o w s   S e r v e r   2 0 1 2  W i n d o w s   8 . 1  W i n d o w s   S e r v e r   2 0 1 2   R 2  W i n 3 2   e r r o r :   % s   ( % u ) % s % s  L i b r a r y   n o t   f o u n d :   % s  F u n c t i o n   n o t   f o u n d :   % s . % s  N o   p a g e   l o a d e d  C a n n o t   r e g i s t e r   a   n i l   p r o v i d e r  I n v a l i d   s e r v i c e   p r o v i d e r   G U I D ) % s   o n l y   s u p p o r t s   s i n k i n g   o f   m e t h o d   c a l l s !   ; D a t a   T L B 1 :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   e n t r i e s E D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   8   e n t r i e s C S h a r e d   2 n d - L e v e l   T L B :   4   K B y t e   p a g e s ,   4 - w a y   a s s o c i a t i v e ,   5 1 2   e n t r i e s D 3 r d - l e v e l   c a c h e :   5 1 2   K B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   1   M B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   2   M B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   1   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   2   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   4   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 3 r d - l e v e l   c a c h e :   1 . 5   M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   3   M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   6   M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   2   M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   4   M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   8   M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 3 r d - l e v e l   c a c h e :   1 2   M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e   Z 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r X 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r C 2 n d - l e v e l   c a c h e :   2   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e A 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e A 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e ? 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e ? 2 n d - l e v e l   c a c h e :   2   M B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e D 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 2 n d - l e v e l   c a c h e :   1   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   1 2 8   e n t r i e s S I n s t r u c t i o n   T L B :   2   M B y t e   p a g e s ,   4 - w a y ,   8   e n t r i e s   o r   4   M B y t e   p a g e s ,   4 - w a y ,   4   e n t r i e s A I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   e n t r i e s ; D a t a   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   1 2 8   e n t r i e s < D a t a   T L B 1 :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   2 5 6   e n t r i e s F D a t a   T L B 0 :   2   M B y t e   o r   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   e n t r i e s / D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   6 4   E n t r i e s 0 D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   1 2 8   E n t r i e s 0 D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   2 5 6   E n t r i e s H 1 s t - l e v e l   d a t a   c a c h e :   1 6   K B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e H 1 s t - l e v e l   d a t a   c a c h e :   8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e I 1 s t - l e v e l   d a t a   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e I 1 s t - l e v e l   d a t a   c a c h e :   3 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e , T r a c e   c a c h e :   1 2   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e , T r a c e   c a c h e :   1 6   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e , T r a c e   c a c h e :   3 2   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e , T r a c e   c a c h e :   6 4   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e : I n s t r u c t i o n   T L B :   2 M / 4 M   p a g e s ,   f u l l y   a s s o c i a t i v e ,   8   e n t r i e s D 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e Z 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r Z 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r   C 3 r d - l e v e l   c a c h e :   8   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   8   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 2 n d - l e v e l   c a c h e :   4   M B y t e s ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   6 M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   8 M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   1 2 M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   1 6 M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 2 n d - l e v e l   c a c h e :   6 M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e * I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   3 2   E n t r i e s A I n s t r u c t i o n   T L B :   4   K B y t e   a n d   2   M B y t e   o r   4   M B y t e   p a g e s ,   6 4   E n t r i e s B I n s t r u c t i o n   T L B :   4   K B y t e   a n d   2   M B y t e   o r   4   M B y t e   p a g e s ,   1 2 8   E n t r i e s B I n s t r u c t i o n   T L B :   4   K B y t e   a n d   2   M B y t e   o r   4   M B y t e   p a g e s ,   2 5 6   E n t r i e s G I n s t r u c t i o n   T L B :   2 - M B y t e   o r   4 - M B y t e   p a g e s ,   f u l l y   a s s o c i a t i v e ,   7   e n t r i e s ; D a t a   T L B 0 :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   1 6   e n t r i e s 7 D a t a   T L B 0 :   4   K B y t e   p a g e s ,   4 - w a y   a s s o c i a t i v e ,   1 6   e n t r i e s 7 D a t a   T L B 0 :   4   K B y t e   p a g e s ,   f u l l y   a s s o c i a t i v e ,   1 6   e n t r i e s W 3 r d   l e v e l   c a c h e :   4   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r I 1 s t   l e v e l   d a t a   c a c h e :   3 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e P 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   3 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   1 9 2   K B y t e s ,   6 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   2 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   3 8 4   K B y t e s ,   6 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e X N o   2 n d - l e v e l   c a c h e   o r ,   i f   p r o c e s s o r   c o n t a i n s   a   v a l i d   2 n d - l e v e l   c a c h e ,   n o   3 r d - l e v e l   c a c h e E 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e C 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e C 2 n d - l e v e l   c a c h e :   2   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   4   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e @ I n s t r u c t i o n   T L B :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   2   e n t r i e s : D a t a   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   e n t r i e s 9 D a t a   T L B :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   8   e n t r i e s ; D a t a   T L B 1 :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   e n t r i e s O 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e P 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e P 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   3 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e H 1 s t   l e v e l   d a t a   c a c h e :   8   K B y t e s ,   2 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e @ I n s t r u c t i o n   T L B :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   4   e n t r i e s I 1 s t   l e v e l   d a t a   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e I 1 s t   l e v e l   d a t a   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e I 1 s t   l e v e l   d a t a   c a c h e :   2 4   K B y t e s ,   6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 2 n d   l e v e l   c a c h e :   2 5 6   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e Y 3 r d   l e v e l   c a c h e :   5 1 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r W 3 r d   l e v e l   c a c h e :   1   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r W 3 r d   l e v e l   c a c h e :   2   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r  P a c k a g e  L i b r a r y 
 N e v e r B u i l d 
 D e s i g n O n l y  R u n O n l y  I g n o r e D u p U n i t s  D e l p h i   3   o r   C + +   B u i l d e r   3 	 U n d e f i n e d  C + +   B u i l d e r   4   o r   l a t e r  D e l p h i   4   o r   l a t e r  M a i n  W e a k  O r g W e a k  I m p l i c i t  N u l l   d e s c r i p t o r A I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   e n t r i e s    N a t i v e  G U I  C o n s o l e  O S / 2  P o s i x 
 R e s e r v e d   8  U N K N O W N  C O F F  C O D E V I E W  F P O  M I S C 	 E X C E P T I O N  F I X U P  O M A P _ T O _ S R C  O M A P _ F R O M _ S R C 
 E x e c u t a b l e    T H U M B  A M 3 3  I B M   P o w e r P C   L i t t l e - E n d i a n  I B M   P o w e r P C   F P  I n t e l   6 4  M I P S 1 6  A L P H A 6 4  M I P S F P U 	 M I P S F P U 1 6  I n f i n e o n  C E F  E F I   B y t e   C o d e 
 A M D 6 4   ( K 8 )  M 3 2 R   l i t t l e - e n d i a n  C E E  U n k n o w n   
 C S D V e r s i o n  R e s e r v e d  E d i t L i s t  U n k n o w n 	 I n t e l   3 8 6  M I P S   l i t t l e - e n d i a n   R 3 0 0 0  M I P S   l i t t l e - e n d i a n   R 4 0 0 0  M I P S   l i t t l e - e n d i a n   R 1 0 0 0 0  M I P S   l i t t l e - e n d i a n   W C E   v 2 	 A l p h a _ A X P  S H 3   l i t t l e - e n d i a n  S H 3   D S P  S H 3 E   l i t t l e - e n d i a n  S H 4   l i t t l e - e n d i a n  S H 5  A R M   L i t t l e - E n d i a n  S i z e   o f   S t a c k   C o m m i t  S i z e   o f   H e a p   R e s e r v e  S i z e   o f   H e a p   C o m m i t  L o a d e r   F l a g s  N u m b e r   o f   R V A  V e r s i o n  G l o b a l F l a g s C l e a r  G l o b a l F l a g s S e t  C r i t i c a l S e c t i o n D e f a u l t T i m e o u t  D e C o m m i t F r e e B l o c k T h r e s h o l d  D e C o m m i t T o t a l F r e e T h r e s h o l d  L o c k P r e f i x T a b l e  M a x i m u m A l l o c a t i o n S i z e  V i r t u a l M e m o r y T h r e s h o l d  P r o c e s s H e a p F l a g s  P r o c e s s A f f i n i t y M a s k    A d d r e s s   o f   E n t r y   P o i n t  B a s e   o f   C o d e  B a s e   o f   D a t a 
 I m a g e   B a s e  S e c t i o n   A l i g n m e n t  F i l e   A l i g n m e n t  O p e r a t i n g   S y s t e m   V e r s i o n  I m a g e   V e r s i o n  S u b s y s t e m   V e r s i o n  W i n 3 2   V e r s i o n  S i z e   o f   I m a g e  S i z e   o f   H e a d e r s  C h e c k S u m 	 S u b s y s t e m  D l l   C h a r a c t e r i s t i c s  S i z e   o f   S t a c k   R e s e r v e    D e l a y   l o a d   i m p o r t  C O M   r u n - t i m e  r e s e r v e d   [ % . 2 d ] 	 S i g n a t u r e  M a c h i n e  N u m b e r   o f   S e c t i o n s  T i m e   D a t e   S t a m p  S y m b o l s   P o i n t e r  N u m b e r   o f   S y m b o l s  S i z e   o f   O p t i o n a l   H e a d e r  C h a r a c t e r i s t i c s  M a g i c  L i n k e r   V e r s i o n  S i z e   o f   C o d e  S i z e   o f   I n i t i a l i z e d   D a t a  S i z e   o f   U n i n i t i a l i z e d   D a t a  N o t   a   r e s o u r c e   d i r e c t o r y , F e a t u r e   i s   n o t   a v a i l a b l e   f o r   a t t a c h e d   i m a g e s  S e c t i o n   " % s "   n o t   f o u n d  E x p o r t s  I m p o r t s 	 R e s o u r c e s 
 E x c e p t i o n s  S e c u r i t y  B a s e   R e l o c a t i o n s  D e b u g  D e s c r i p t i o n  M a c h i n e   V a l u e  T L S  L o a d   c o n f i g u r a t i o n  B o u n d   I m p o r t  I A T % T h i s   w i n d o w s   v e r s i o n   i s   n o t   s u p p o r t e d & T h e   w i n d o w   w i t h   h a n d l e   % d   i s   n o t   v a l i d # T h e   p r o c e s s   w i t h   I D   % d   i s   n o t   v a l i d & T h e   M o d u l e   w i t h   h a n d l e   % d   i s   n o t   v a l i d $ F i l e   c o n t a i n s   n o   v e r s i o n   i n f o r m a t i o n  T h e   f i l e   % s   d o e s   n o t   e x i s t  I l l e g a l   l a n g u a g e   i n d e x  N o   v a l u e   w a s   s u p p l i e d  T h e   v a l u e   % s   w a s   n o t   f o u n d .  F a i l e d   t o   c r e a t e   F i l e M a p p i n g   F a i l e d   t o   c r e a t e   F i l e M a p p i n g V i e w  F a i l e d   t o   o b t a i n   s i z e   o f   f i l e  S t r e a m   i s   r e a d - o n l y  C a n n o t   o p e n   f i l e   " % s "  T h i s   i s   n o t   a   P E   f o r m a t  U n k n o w n   P E   t a r g e t    T h e r e   i s   n o   s u c h   p a l e t t e   e n t r y . d T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   a n   u n k n o w n   c r i t i c a l   p a r t   w h i c h   c o u l d   n o t   b e   d e c o d e d . p T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   e n c o d e d   w i t h   a n   u n k n o w n   c o m p r e s s i o n   s c h e m e   w h i c h   c o u l d   n o t   b e   d e c o d e d . c T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   u s e s   a n   u n k n o w n   i n t e r l a c e   s c h e m e   w h i c h   c o u l d   n o t   b e   d e c o d e d . - T h e   c h u n k s   m u s t   b e   c o m p a t i b l e   t o   b e   a s s i g n e d . j T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   i n v a l i d   b e c a u s e   t h e   d e c o d e r   f o u n d   a n   u n e x p e c t e d   e n d   o f   t h e   f i l e . 8 T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   n o   d a t a . ] T h e   p r o g r a m   t r i e d   t o   a d d   a   e x i s t e n t   c r i t i c a l   c h u n k   t o   t h e   c u r r e n t   i m a g e   w h i c h   i s   n o t   a l l o w e d . I I t ' s   n o t   a l l o w e d   t o   a d d   a   n e w   c h u n k   b e c a u s e   t h e   c u r r e n t   i m a g e   i s   i n v a l i d . 7 T h e   p n g   i m a g e   c o u l d   n o t   b e   l o a d e d   f r o m   t h e   r e s o u r c e   I D . o S o m e   o p e r a t i o n   c o u l d   n o t   b e   p e r f o r m e d   b e c a u s e   t h e   s y s t e m   i s   o u t   o f   r e s o u r c e s .   C l o s e   s o m e   w i n d o w s   a n d   t r y   a g a i n . � S e t t i n g   b i t   t r a n s p a r e n c y   c o l o r   i s   n o t   a l l o w e d   f o r   p n g   i m a g e s   c o n t a i n i n g   a l p h a   v a l u e   f o r   e a c h   p i x e l   ( C O L O R _ R G B A L P H A   a n d   C O L O R _ G R A Y S C A L E A L P H A ) O T h i s   o p e r a t i o n   i s   n o t   v a l i d   b e c a u s e   t h e   c u r r e n t   i m a g e   c o n t a i n s   n o   v a l i d   h e a d e r . 4 T h e   n e w   s i z e   p r o v i d e d   f o r   i m a g e   r e s i z i n g   i s   i n v a l i d . o T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   i n v a l i d   i m a g e   t y p e   p a r a m e t e r s   h a v e   b e i n g   p r o v i d e d . ( F a i l e d   t o   g e t   A N S I   r e p l a c e m e n t   c h a r a c t e r   + M i s m a t c h e d   p a r a m a t e r s   t o   R e g i s t e r C h i l d N o d e s 0 E l e m e n t   " % s "   d o e s   n o t   c o n t a i n   a   s i n g l e   t e x t   n o d e 4 D O M   I m p l e m e n t a t i o n   d o e s   n o t   s u p p o r t   I D O M P a r s e O p t i o n s # I t e m T a g   p r o p e r t y   i s   n o t   i n i t i a l i z e d  N o d e   i s   r e a d o n l y C R e f r e s h   i s   o n l y   s u p p o r t e d   i f   t h e   F i l e N a m e   o r   X M L   p r o p e r t i e s   a r e   s e t  F i l e N a m e   c a n n o t   b e   b l a n k  L i n e j T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   v a l i d   b e c a u s e   i t   c o n t a i n s   i n v a l i d   p i e c e s   o f   d a t a   ( c r c   e r r o r ) y T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o u l d   n o t   b e   l o a d e d   b e c a u s e   o n e   o f   i t s   m a i n   p i e c e   o f   d a t a   ( i h d r )   m i g h t   b e   c o r r u p t e d U T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   i n v a l i d   b e c a u s e   i t   h a s   m i s s i n g   i m a g e   p a r t s . [ C o u l d   n o t   d e c o m p r e s s   t h e   i m a g e   b e c a u s e   i t   c o n t a i n s   i n v a l i d   c o m p r e s s e d   d a t a .  
   D e s c r i p t i o n :   B T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   a n   i n v a l i d   p a l e t t e . � T h e   f i l e   b e i n g   r e a d   i s   n o t   a   v a l i d   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   b e c a u s e   i t   c o n t a i n s   a n   i n v a l i d   h e a d e r .   T h i s   f i l e   m a y   b e   c o r r u p t e d ,   t r y   o b t a i n i n g   i t   a g a i n n T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   s u p p o r t e d   o r   i t   m i g h t   b e   i n v a l i d .  
 ( I H D R   c h u n k   i s   n o t   t h e   f i r s t ) � T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   s u p p o r t e d   b e c a u s e   e i t h e r   i t s   w i d t h   o r   h e i g h t   e x c e e d s   t h e   m a x i m u m   s i z e   o f   6 5 5 3 5   p i x e l s .  M o r e   B u t t o n s | J A   T T B D o c k   c o n t r o l   c a n n o t   b e   p l a c e d   i n s i d e   a   t o o l   w i n d o w   o r   a n o t h e r   T T B D o c k C C a n n o t   c h a n g e   P o s i t i o n   o f   a   T T B D o c k   i f   i t   a l r e a d y   c o n t a i n s   c o n t r o l s G C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   N a m e   p r o p e r t y   i s   n o t   s e t O C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   D o c k e d T o ' s   N a m e   p r o p e r t y   n o t   s e t ) " % s "   D O M I m p l e m e n t a t i o n   a l r e a d y   r e g i s t e r e d  N o   m a t c h i n g   D O M   V e n d o r :   " % s " < S e l e c t e d   D O M   V e n d o r   d o e s   n o t   s u p p o r t   t h i s   p r o p e r t y   o r   m e t h o d ; P r o p e r t y   o r   M e t h o d   " % s "   i s   n o t   s u p p o r t e d   b y   D O M   V e n d o r   " % s "  N o d e   c a n n o t   b e   n u l l   M i c r o s o f t   M S X M L   i s   n o t   i n s t a l l e d  N o   a c t i v e   d o c u m e n t  N o d e   " % s "   n o t   f o u n d  I D O M N o d e   r e q u i r e d . A t t r i b u t e s   a r e   n o t   s u p p o r t e d   o n   t h i s   n o d e   t y p e  I n v a l i d   n o d e   t y p e  � n d r a d  A t t r  E x t  % s   � r   e n   o g i l t i g   e n h e t s b o k s t a v .  R � t t i g h e t e r  � g a r e  G r u p p  M � l   l � n k  F i l t y p  & K o p i e r a   h i t  & F l y t t a   h i t  & S k a p a   g e n v � g   h i t  & A v b r y t  T o o l b a r   i t e m   i n d e x   o u t   o f   r a n g e  T o o l b a r   i t e m   a l r e a d y   i n s e r t e d ? A n   i t e m   v i e w e r   a s s o c i a t e d   t h e   s p e c i f i e d   i t e m   c o u l d   n o t   b e   f o u n d    M B  G B ) K a n   i n t e   b y t a   n a m n   p �   f i l   e l l e r   k a t a l o g :    F i l e n   f i n n s   r e d a n :   % F i l n a m n e t   i n n e h � l l e r   o g i l t i g a   t e c k e n :  F i l   % s  % u   F i l e r  % u   K a t a l o g e r  H u v u d k a t a l o g  D r a g D r o p   E r r o r :   % d  E n h e t   ' % s : '   � r   i n t e   k l a r .  K a t a l o g e n   ' % s '   f i n n s   i n t e .  /   < r o o t >  N a m n  S t o r l e k  F i l t y p    U n a b l e   t o   c r e a t e   d i r e c t o r y  I n v a l i d   s o u r c e   a r r a y  I n v a l i d   d e s t i n a t i o n   a r r a y " C h a r a c t e r   i n d e x   o u t   o f   b o u n d s   ( % d )  S t a r t   i n d e x   o u t   o f   b o u n d s   ( % d )  I n v a l i d   c o u n t   ( % d )  I n v a l i d   d e s t i n a t i o n   i n d e x   ( % d )  I n v a l i d   c o d e   p a g e  I n v a l i d   e n c o d i n g   n a m e N N o   m a p p i n g   f o r   t h e   U n i c o d e   c h a r a c t e r   e x i s t s   i n   t h e   t a r g e t   m u l t i - b y t e   c o d e   p a g e  B l � d d r a  A l l a   f i l e r   ( * . * ) | * . *  O g i l t i g t   f i l n a m n   -   % s # K a n   i n t e   h i t t a   n � g o n   g i l t i g   s � k v � g .  B  K B    N o v e m b e r  D e c e m b e r  S u n  M o n  T u e  W e d  T h u  F r i  S a t  S u n d a y  M o n d a y  T u e s d a y 	 W e d n e s d a y  T h u r s d a y  F r i d a y  S a t u r d a y    J u l  A u g  S e p  O c t  N o v  D e c  J a n u a r y  F e b r u a r y  M a r c h  A p r i l  M a y  J u n e  J u l y  A u g u s t 	 S e p t e m b e r  O c t o b e r ( M o n i t o r   s u p p o r t   f u n c t i o n   n o t   i n i t i a l i z e d  F e a t u r e   n o t   i m p l e m e n t e d   M e t h o d   c a l l e d   o n   d i s p o s e d   o b j e c t  % s   ( % s ,   l i n e   % d )  A b s t r a c t   E r r o r ? A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p   i n   m o d u l e   ' % s ' .   % s   o f   a d d r e s s   % p 2 C a n n o t   a c c e s s   p a c k a g e   i n f o r m a t i o n   f o r   p a c k a g e   ' % s '  C a n ' t   l o a d   p a c k a g e   % s .  
 % s  S y s t e m f e l .   K o d :   % d .  
 % s % s * E t t   a n r o p   t i l l   e n   O S   f u n k t i o n   m i s s l y c k a d e s  J a n  F e b  M a r  A p r  M a y  J u n   , C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   i s   o u t   o f   r a n g e / C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   a l r e a d y   u s e d   b y   % s * C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   i s   n o t   u s a b l e 2 T o o   m a n y   c u s t o m   v a r i a n t   t y p e s   h a v e   b e e n   r e g i s t e r e d 5 C o u l d   n o t   c o n v e r t   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s ) = O v e r f l o w   w h i l e   c o n v e r t i n g   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s )  V a r i a n t   o v e r f l o w  I n v a l i d   a r g u m e n t  I n v a l i d   v a r i a n t   t y p e  O p e r a t i o n   n o t   s u p p o r t e d  U n e x p e c t e d   v a r i a n t   e r r o r  E x t e r n a l   e x c e p t i o n   % x  A s s e r t i o n   f a i l e d  I n t e r f a c e   n o t   s u p p o r t e d  E x c e p t i o n   i n   s a f e c a l l   m e t h o d  O b j e c t   l o c k   n o t   o w n e d    A p p l i c a t i o n   E r r o r 1 F o r m a t   ' % s '   i n v a l i d   o r   i n c o m p a t i b l e   w i t h   a r g u m e n t  N o   a r g u m e n t   f o r   f o r m a t   ' % s ' " V a r i a n t   m e t h o d   c a l l s   n o t   s u p p o r t e d  R e a d  W r i t e 	 E x e c u t i o n  I n v a l i d   a c c e s s  F o r m a t   s t r i n g   t o o   l o n g $ E r r o r   c r e a t i n g   v a r i a n t   o r   s a f e   a r r a y ) V a r i a n t   o r   s a f e   a r r a y   i n d e x   o u t   o f   b o u n d s  V a r i a n t   o r   s a f e   a r r a y   i s   l o c k e d  I n v a l i d   v a r i a n t   t y p e   c o n v e r s i o n  I n v a l i d   v a r i a n t   o p e r a t i o n  I n v a l i d   N U L L   v a r i a n t   o p e r a t i o n % I n v a l i d   v a r i a n t   o p e r a t i o n   ( % s % . 8 x ) 
 % s  D i v i s i o n   b y   z e r o  R a n g e   c h e c k   e r r o r  I n t e g e r   o v e r f l o w   I n v a l i d   f l o a t i n g   p o i n t   o p e r a t i o n  F l o a t i n g   p o i n t   d i v i s i o n   b y   z e r o  F l o a t i n g   p o i n t   o v e r f l o w  F l o a t i n g   p o i n t   u n d e r f l o w  I n v a l i d   p o i n t e r   o p e r a t i o n  I n v a l i d   c l a s s   t y p e c a s t 0 A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p .   % s   o f   a d d r e s s   % p  A c c e s s   v i o l a t i o n  S t a c k   o v e r f l o w  C o n t r o l - C   h i t  P r i v i l e g e d   i n s t r u c t i o n  O p e r a t i o n   a b o r t e d ( E x c e p t i o n   % s   i n   m o d u l e   % s   a t   % p .  
 % s % s  
 ! ' % s '   i s   n o t   a   v a l i d   i n t e g e r   v a l u e ( ' % s '   i s   n o t   a   v a l i d   f l o a t i n g   p o i n t   v a l u e  ' % s '   � r   i n g e t   g i l t i g t   d a t u m  ' % s '   � r   i n g e n   g i l t i g   t i d # ' % s '   � r   i n g e t   g i l t i g t   d a t u m   o c h   t i d   ' % d . % d '   i s   n o t   a   v a l i d   t i m e s t a m p  ' % s '   i s   n o t   a   v a l i d   G U I D   v a l u e  I n v a l i d   a r g u m e n t   t o   t i m e   e n c o d e  I n v a l i d   a r g u m e n t   t o   d a t e   e n c o d e  O u t   o f   m e m o r y  I / O   e r r o r   % d  T o o   m a n y   o p e n   f i l e s  F i l e   a c c e s s   d e n i e d  R e a d   b e y o n d   e n d   o f   f i l e 	 D i s k   f u l l  I n v a l i d   n u m e r i c   i n p u t  W i n d o w s   S e r v e r   2 0 0 3   R 2  W i n d o w s   S e r v e r   2 0 1 2  W i n d o w s   S e r v e r   2 0 1 2   R 2 	 W i n d o w s   8  W i n d o w s   8 . 1  O b s e r v e r   i s   n o t   s u p p o r t e d L C a n n o t   h a v e   m u l t i p l e   s i n g l e   c a s t   o b s e r v e r s   a d d e d   t o   t h e   o b s e r v e r s   c o l l e c t i o n 4 T h e   o b j e c t   d o e s   n o t   i m p l e m e n t   t h e   o b s e r v e r   i n t e r f a c e G N o   s i n g l e   c a s t   o b s e r v e r   w i t h   I D   % d   w a s   a d d e d   t o   t h e   o b s e r v e r   c o l l e c t i o n F N o   m u l t i   c a s t   o b s e r v e r   w i t h   I D   % d   w a s   a d d e d   t o   t h e   o b s e r v e r   c o l l e c t i o n  O b s e r v e r   i s   n o t   a v a i l a b l e  T h e   l o c a t i o n   s e n s o r   i s   s t a r t e d  I n v a l i d   d a t e   s t r i n g :   % s  I n v a l i d   t i m e   s t r i n g :   % s  I n v a l i d   t i m e   O f f s e t   s t r i n g :   % s 	 < u n k n o w n >    P a r a m e t e r   c o u n t   m i s m a t c h < T y p e   ' % s '   i s   n o t   d e c l a r e d   i n   t h e   i n t e r f a c e   s e c t i o n   o f   a   u n i t 7 V A R   a n d   O U T   a r g u m e n t s   m u s t   m a t c h   p a r a m e t e r   t y p e   e x a c t l y , S p e c i f i e d   L o g i n   C r e d e n t i a l   S e r v i c e   n o t   f o u n d " % s   ( V e r s i o n   % d . % d ,   B u i l d   % d ,   % 5 : s ) : % s   S e r v i c e   P a c k   % 4 : d   ( V e r s i o n   % 1 : d . % 2 : d ,   B u i l d   % 3 : d ,   % 5 : s )  3 2 - b i t   E d i t i o n  6 4 - b i t   E d i t i o n  W i n d o w s  W i n d o w s   V i s t a  W i n d o w s   S e r v e r   2 0 0 8 	 W i n d o w s   7  W i n d o w s   S e r v e r   2 0 0 8   R 2  W i n d o w s   2 0 0 0 
 W i n d o w s   X P  W i n d o w s   S e r v e r   2 0 0 3 b T h e   d u r a t i o n   c a n n o t   b e   r e t u r n e d   b e c a u s e   t h e   a b s o l u t e   v a l u e   e x c e e d s   t h e   v a l u e   o f   T T i m e S p a n . M a x V a l u e  V a l u e   c a n n o t   b e   N a N 3 N e g a t i n g   t h e   m i n i m u m   v a l u e   o f   a   T i m e s p a n   i s   i n v a l i d  I n v a l i d   T i m e s p a n   f o r m a t  T i m e s p a n   e l e m e n t   t o o   l o n g # N o   c o n t e x t - s e n s i t i v e   h e l p   i n s t a l l e d  N o   h e l p   f o u n d   f o r   c o n t e x t   % d  U n a b l e   t o   o p e n   I n d e x  U n a b l e   t o   o p e n   S e a r c h " U n a b l e   t o   f i n d   a   T a b l e   o f   C o n t e n t s $ N o   t o p i c - b a s e d   h e l p   s y s t e m   i n s t a l l e d  N o   h e l p   f o u n d   f o r   % s  A r g u m e n t   o u t   o f   r a n g e  I t e m   n o t   f o u n d  D u p l i c a t e s   n o t   a l l o w e d 5 I n s u f f i c i e n t   R T T I   a v a i l a b l e   t o   s u p p o r t   t h i s   o p e r a t i o n  T h e   s p e c i f i e d   p a t h   i s   t o o   l o n g   T h e   s p e c i f i e d   p a t h   w a s   n o t   f o u n d   T h e   p a t h   f o r m a t   i s   n o t   s u p p o r t e d  T h e   d r i v e   c a n n o t   b e   f o u n d   T h e   s p e c i f i e d   f i l e   w a s   n o t   f o u n d ! T h e   s p e c i f i e d   f i l e   a l r e a d y   e x i s t s  ? W T h e   g i v e n   " % s "   l o c a l   t i m e   i s   i n v a l i d   ( s i t u a t e d   w i t h i n   t h e   m i s s i n g   p e r i o d   p r i o r   t o   D S T ) . $ N o   h e l p   v i e w e r   t h a t   s u p p o r t s   f i l t e r s 8 S t r i n g   i n d e x   o u t   o f   r a n g e   ( % d ) .     M u s t   b e   > =   % d   a n d   < =   % d \ I n v a l i d   U T F 3 2   c h a r a c t e r   v a l u e .     M u s t   b e   > =   0   a n d   < =   $ 1 0 F F F F ,   e x c l u d i n g   s u r r o g a t e   p a i r   r a n g e s r H i g h   s u r r o g a t e   c h a r   w i t h o u t   a   f o l l o w i n g   l o w   s u r r o g a t e   c h a r   a t   i n d e x :   % d .   C h e c k   t h a t   t h e   s t r i n g   i s   e n c o d e d   p r o p e r l y r L o w   s u r r o g a t e   c h a r   w i t h o u t   a   p r e c e d i n g   h i g h   s u r r o g a t e   c h a r   a t   i n d e x :   % d .   C h e c k   t h a t   t h e   s t r i n g   i s   e n c o d e d   p r o p e r l y 2 L e n g t h   o f   S t r i n g s   a n d   O b j e c t s   a r r a y s   m u s t   b e   e q u a l  I n v a l i d   T i m e o u t   v a l u e :   % s  T i m e s p a n   t o o   l o n g  S t r i n g   e x p e c t e d  % s   e x p e c t e d $ % s   n o t   i n   a   c l a s s   r e g i s t r a t i o n   g r o u p  P r o p e r t y   % s   d o e s   n o t   e x i s t  S t r e a m   w r i t e   e r r o r  T h r e a d   c r e a t i o n   e r r o r :   % s  T h r e a d   E r r o r :   % s   ( % d ) - C a n n o t   t e r m i n a t e   a n   e x t e r n a l l y   c r e a t e d   t h r e a d , C a n n o t   w a i t   f o r   a n   e x t e r n a l l y   c r e a t e d   t h r e a d 2 C a n n o t   c a l l   S t a r t   o n   a   r u n n i n g   o r   s u s p e n d e d   t h r e a d ; C a n n o t   c a l l   C h e c k T e r m i n a t e d   o n   a n   e x t e r n a l l y   c r e a t e d   t h r e a d 9 C a n n o t   c a l l   S e t R e t u r n V a l u e   o n   a n   e x t e r n a l l y   c r e a t e   t h r e a d  P a r a m e t e r   % s   c a n n o t   b e   n i l ' P a r a m e t e r   % s   c a n n o t   b e   a   n e g a t i v e   v a l u e * I n p u t   b u f f e r   e x c e e d e d   f o r   % s   =   % d ,   % s   =   % d  I n v a l i d   c h a r a c t e r s   i n   p a t h  L i s t   i n d e x   o u t   o f   b o u n d s   ( % d ) + O u t   o f   m e m o r y   w h i l e   e x p a n d i n g   m e m o r y   s t r e a m ) % s   h a s   n o t   b e e n   r e g i s t e r e d   a s   a   C O M   c l a s s  N u m b e r   e x p e c t e d  A N S I   o r   U T F 8   e n c o d i n g   e x p e c t e d  % s   o n   l i n e   % d  E r r o r   r e a d i n g   % s % s % s :   % s  S t r e a m   r e a d   e r r o r  P r o p e r t y   i s   r e a d - o n l y  F a i l e d   t o   c r e a t e   k e y   % s  F a i l e d   t o   g e t   d a t a   f o r   ' % s '  I n v a l i d   c o m p o n e n t   r e g i s t r a t i o n  F a i l e d   t o   s e t   d a t a   f o r   ' % s '  R e s o u r c e   % s   n o t   f o u n d  % s . S e e k   n o t   i m p l e m e n t e d $ O p e r a t i o n   n o t   a l l o w e d   o n   s o r t e d   l i s t  U n a b l e   t o   w r i t e   t o   % s  I n v a l i d   b i n a r y   v a l u e  I n v a l i d   f i l e   n a m e   -   % s  I n v a l i d   s t r e a m   f o r m a t  ' % s '   i s   a n   i n v a l i d   m a s k   a t   ( % d ) $ ' ' % s ' '   i s   n o t   a   v a l i d   c o m p o n e n t   n a m e  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   p r o p e r t y   e l e m e n t :   % s  I n v a l i d   p r o p e r t y   p a t h  I n v a l i d   p r o p e r t y   t y p e :   % s  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   d a t a   t y p e   f o r   ' % s '  I n v a l i d   s t r i n g   c o n s t a n t  L i n e   t o o   l o n g   L i s t   c a p a c i t y   o u t   o f   b o u n d s   ( % d )  L i s t   c o u n t   o u t   o f   b o u n d s   ( % d ) 7 D i s p a t c h   m e t h o d s   d o   n o t   s u p p o r t   m o r e   t h a n   6 4   p a r a m e t e r s  D C O M   n o t   i n s t a l l e d  A n c e s t o r   f o r   ' % s '   n o t   f o u n d  C a n n o t   a s s i g n   a   % s   t o   a   % s  B i t s   i n d e x   o u t   o f   r a n g e * C a n ' t   w r i t e   t o   a   r e a d - o n l y   r e s o u r c e   s t r e a m  ' ' % s ' '   e x p e c t e d E C h e c k S y n c h r o n i z e   c a l l e d   f r o m   t h r e a d   $ % x ,   w h i c h   i s   N O T   t h e   m a i n   t h r e a d  C l a s s   % s   n o t   f o u n d  A   c l a s s   n a m e d   % s   a l r e a d y   e x i s t s % L i s t   d o e s   n o t   a l l o w   d u p l i c a t e s   ( $ 0 % x ) # A   c o m p o n e n t   n a m e d   % s   a l r e a d y   e x i s t s % S t r i n g   l i s t   d o e s   n o t   a l l o w   d u p l i c a t e s  C a n n o t   c r e a t e   f i l e   " % s " .   % s  C a n n o t   o p e n   f i l e   " % s " .   % s  I d e n t i f i e r   e x p e c t e d 4 Y o u   m u s t   b e   i n   S h o w C h e c k b o x   m o d e   t o   s e t   t o   t h i s   d a t e # F a i l e d   t o   s e t   c a l e n d a r   d a t e   o r   t i m e % F a i l e d   t o   s e t   m a x i m u m   s e l e c t i o n   r a n g e $ F a i l e d   t o   s e t   c a l e n d a r   m i n / m a x   r a n g e % F a i l e d   t o   s e t   c a l e n d a r   s e l e c t e d   r a n g e 3 A   r e g u l a r   e x p r e s s i o n   s p e c i f i e d   i n   R e g E x   i s   r e q u i r e d , E r r o r   i n   r e g u l a r   e x p r e s s i o n   a t   o f f s e t   % d :   % s  E r r o r   s t u d y i n g   t h e   r e g e x :   % s  S u c c e s s f u l   m a t c h   r e q u i r e d  S t r i n g s   p a r a m e t e r   c a n n o t   b e   n i l  I n v a l i d   i n d e x   t y p e  I n d e x   o u t   o f   b o u n d s   ( % d )  I n v a l i d   g r o u p   n a m e   ( % s )  O L E   e r r o r   % . 8 x . M e t h o d   ' % s '   n o t   s u p p o r t e d   b y   a u t o m a t i o n   o b j e c t / V a r i a n t   d o e s   n o t   r e f e r e n c e   a n   a u t o m a t i o n   o b j e c t " F a i l e d   t o   s e t   t a b   " % s "   a t   i n d e x   % d   F a i l e d   t o   s e t   o b j e c t   a t   i n d e x   % d < M u l t i L i n e   m u s t   b e   T r u e   w h e n   T a b P o s i t i o n   i s   t p L e f t   o r   t p R i g h t  I n v a l i d   i t e m   l e v e l   a s s i g n m e n t   I n v a l i d   l e v e l   ( % d )   f o r   i t e m   " % s "  I n v a l i d   i n d e x  U n a b l e   t o   i n s e r t   a n   i t e m  I n v a l i d   o w n e r  R i c h E d i t   l i n e   i n s e r t i o n   e r r o r  F a i l e d   t o   L o a d   S t r e a m  F a i l e d   t o   S a v e   S t r e a m   % s   i s   a l r e a d y   a s s o c i a t e d   w i t h   % s E % d   i s   a n   i n v a l i d   P a g e I n d e x   v a l u e .     P a g e I n d e x   m u s t   b e   b e t w e e n   0   a n d   % d = T h i s   c o n t r o l   r e q u i r e s   v e r s i o n   4 . 7 0   o r   g r e a t e r   o f   C O M C T L 3 2 . D L L  D a t e   e x c e e d s   m a x i m u m   o f   % s  D a t e   i s   l e s s   t h a n   m i n i m u m   o f   % s    % s   p a r a m e t e r   c a n n o t   b e   n i l 0 A   S t y l e H o o k   c l a s s   h a s   n o t   b e e n   r e g i s t e r e d   f o r   % s # F e a t u r e   n o t   s u p p o r t e d   b y   t h i s   s t y l e  S t y l e   ' % s '   i s   n o t   r e g i s t e r e d " C a n n o t   u n r e g i s t e r   t h e   s y s t e m   s t y l e  S t y l e   n o t   r e g i s t e r e d " ' % s '   i s   n o t   a   v a l i d   p r o p e r t y   v a l u e  O L E   c o n t r o l   a c t i v a t i o n   f a i l e d * C o u l d   n o t   o b t a i n   O L E   c o n t r o l   w i n d o w   h a n d l e % L i c e n s e   i n f o r m a t i o n   f o r   % s   i s   i n v a l i d P L i c e n s e   i n f o r m a t i o n   f o r   % s   n o t   f o u n d .   Y o u   c a n n o t   u s e   t h i s   c o n t r o l   i n   d e s i g n   m o d e N U n a b l e   t o   r e t r i e v e   a   p o i n t e r   t o   a   r u n n i n g   o b j e c t   r e g i s t e r e d   w i t h   O L E   f o r   % s / % s  F a i l e d   t o   c l e a r   t a b   c o n t r o l   F a i l e d   t o   d e l e t e   t a b   a t   i n d e x   % d " F a i l e d   t o   r e t r i e v e   t a b   a t   i n d e x   % d   F a i l e d   t o   g e t   o b j e c t   a t   i n d e x   % d  R a d i o B u t t o n % d  C a p t i o n   c a n n o t   b e   e m p t y : C a t e g o r y P a n e l   m u s t   h a v e   a   C a t e g o r y P a n e l G r o u p   a s   i t s   p a r e n t = O n l y   C a t e g o r y P a n e l s   c a n   b e   i n s e r t e d   i n t o   a   C a t e g o r y P a n e l G r o u p  N o   h e l p   k e y w o r d   s p e c i f i e d .  U n a b l e   t o   l o a d   s t y l e   ' % s '  U n a b l e   t o   l o a d   s t y l e s :   % s  S t y l e   ' % s '   a l r e a d y   r e g i s t e r e d # S t y l e   c l a s s   ' % s '   a l r e a d y   r e g i s t e r e d  S t y l e   ' % s '   n o t   f o u n d  S t y l e   c l a s s   ' % s '   n o t   f o u n d  I n v a l i d   s t y l e   h a n d l e  I n v a l i d   s t y l e   f o r m a t  V C L   S t y l e   F i l e ) C l a s s   ' % s '   i s   a l r e a d y   r e g i s t e r e d   f o r   ' % s ' % C l a s s   ' % s '   i s   n o t   r e g i s t e r e d   f o r   ' % s '    L o g i n 	 S e p a r a t o r  E r r o r   s e t t i n g   % s . C o u n t 8 L i s t b o x   ( % s )   s t y l e   m u s t   b e   v i r t u a l   i n   o r d e r   t o   s e t   C o u n t # N o   O n G e t I t e m   e v e n t   h a n d l e r   a s s i g n e d  " % s "   i s   a n   i n v a l i d   p a t h  A N S I  A S C I I  U n i c o d e  B i g   E n d i a n   U n i c o d e  U T F - 8  U T F - 7 % C a n n o t   r e m o v e   s h e l l   n o t i f i c a t i o n   i c o n " P a g e C o n t r o l   m u s t   f i r s t   b e   a s s i g n e d " % s   r e q u i r e s   W i n d o w s   V i s t a   o r   l a t e r  B u t t o n % d   . T h e r e   i s   n o   d e f a u l t   p r i n t e r   c u r r e n t l y   s e l e c t e d / M e n u   ' % s '   i s   a l r e a d y   b e i n g   u s e d   b y   a n o t h e r   f o r m  P i c t u r e :    ( % d x % d )  P r e v i e w  D o c k e d   c o n t r o l   m u s t   h a v e   a   n a m e % E r r o r   r e m o v i n g   c o n t r o l   f r o m   d o c k   t r e e    -   D o c k   z o n e   n o t   f o u n d    -   D o c k   z o n e   h a s   n o   c o n t r o l L E r r o r   l o a d i n g   d o c k   z o n e   f r o m   t h e   s t r e a m .   E x p e c t i n g   v e r s i o n   % d ,   b u t   f o u n d   % d . , M u l t i s e l e c t   m o d e   m u s t   b e   o n   f o r   t h i s   f e a t u r e 7 L e n g t h   o f   v a l u e   a r r a y   m u s t   b e   > =   l e n g t h   o f   p r o m p t   a r r a y  P r o m p t   a r r a y   m u s t   n o t   b e   e m p t y 	 & U s e r n a m e 	 & P a s s w o r d  & D o m a i n    R i g h t  D o w n  I n s  D e l  S h i f t +  C t r l +  A l t +  ( N o n e )  V a l u e   m u s t   b e   b e t w e e n   % d   a n d   % d  A l l  U n a b l e   t o   i n s e r t   a   l i n e  I n v a l i d   c l i p b o a r d   f o r m a t   C l i p b o a r d   d o e s   n o t   s u p p o r t   I c o n s  C a n n o t   o p e n   c l i p b o a r d :   % s  T e x t   e x c e e d s   m e m o   c a p a c i t y + O p e r a t i o n   n o t   s u p p o r t e d   o n   s e l e c t e d   p r i n t e r   	 & I g n o r e r a  & A l l a  N & e j   t i l l   a l l a  J & a   t i l l   a l l a  & S t � n g  B k S p  T a b  E s c  E n t e r  S p a c e  P g U p  P g D n  E n d  H o m e  L e f t  U p 1 F i x e d   c o l u m n   c o u n t   m u s t   b e   l e s s   t h a n   c o l u m n   c o u n t + F i x e d   r o w   c o u n t   m u s t   b e   l e s s   t h a n   r o w   c o u n t & C a n n o t   i n s e r t   o r   d e l e t e   r o w s   f r o m   g r i d  O g i l t i g t   i n p u t v � r d e 9 O g i l t i g t   i n p u t v � r d e .   A n v � n d   E S C   f � r   a t t   a v b r y t a   � n d r i n g a r  V a r n i n g  F e l  I n f o r m a t i o n  B e k r � f t a  & J a  & N e j  O K  A v b r y t  & H j � l p  & A v b r y t  & F � r s � k   i g e n    & N o  & H e l p  & C l o s e  & I g n o r e  & R e t r y  A b o r t  & A l l  C a n n o t   d r a g   a   f o r m 	 M e t a f i l e s  E n h a n c e d   M e t a f i l e s  I c o n s  B i t m a p s  T I F F   I m a g e s  G r i d   t o o   l a r g e   f o r   o p e r a t i o n   T o o   m a n y   r o w s   o r   c o l u m n s   d e l e t e d  G r i d   i n d e x   o u t   o f   r a n g e    M e n u   i n d e x   o u t   o f   r a n g e  M e n u   i n s e r t e d   t w i c e  S u b - m e n u   i s   n o t   i n   m e n u  N o t   e n o u g h   t i m e r s   a v a i l a b l e ! P r i n t e r   i s   n o t   c u r r e n t l y   p r i n t i n g  P r i n t i n g   i n   p r o g r e s s  P r i n t e r   i n d e x   o u t   o f   r a n g e  P r i n t e r   s e l e c t e d   i s   n o t   v a l i d  % s   o n   % s @ G r o u p I n d e x   c a n n o t   b e   l e s s   t h a n   a   p r e v i o u s   m e n u   i t e m ' s   G r o u p I n d e x 5 C a n n o t   c r e a t e   f o r m .   N o   M D I   f o r m s   a r e   c u r r e n t l y   a c t i v e 0 C a n   o n l y   m o d i f y   a n   i m a g e   i f   i t   c o n t a i n s   a   b i t m a p * A   c o n t r o l   c a n n o t   h a v e   i t s e l f   a s   i t s   p a r e n t  O K  A v b r y t  & Y e s    I n v a l i d   i m a g e   s i z e  I n v a l i d   I m a g e L i s t  U n a b l e   t o   R e p l a c e   I m a g e  I n v a l i d   I m a g e L i s t   I n d e x ) F a i l e d   t o   r e a d   I m a g e L i s t   d a t a   f r o m   s t r e a m ( F a i l e d   t o   w r i t e   I m a g e L i s t   d a t a   t o   s t r e a m $ E r r o r   c r e a t i n g   w i n d o w   d e v i c e   c o n t e x t  E r r o r   c r e a t i n g   w i n d o w   c l a s s + C a n n o t   f o c u s   a   d i s a b l e d   o r   i n v i s i b l e   w i n d o w ! C o n t r o l   ' % s '   h a s   n o   p a r e n t   w i n d o w $ P a r e n t   g i v e n   i s   n o t   a   p a r e n t   o f   ' % s '  C a n n o t   h i d e   a n   M D I   C h i l d   F o r m ) C a n n o t   c h a n g e   V i s i b l e   i n   O n S h o w   o r   O n H i d e " C a n n o t   m a k e   a   v i s i b l e   w i n d o w   m o d a l  S c r o l l b a r   p r o p e r t y   o u t   o f   r a n g e  % s   p r o p e r t y   o u t   o f   r a n g e 0 T a b   p o s i t i o n   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   s t y l e 0 T a b   s t y l e   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   p o s i t i o n  B i t m a p   i m a g e   i s   n o t   v a l i d  I c o n   i m a g e   i s   n o t   v a l i d  M e t a f i l e   i s   n o t   v a l i d  I n v a l i d   p i x e l   f o r m a t  I n v a l i d   i m a g e  S c a n   l i n e   i n d e x   o u t   o f   r a n g e ! C a n n o t   c h a n g e   t h e   s i z e   o f   a n   i c o n % C a n n o t   c h a n g e   t h e   s i z e   o f   a   W I C   I m a g e   I n v a l i d   o p e r a t i o n   o n   T O l e G r a p h i c $ U n k n o w n   p i c t u r e   f i l e   e x t e n s i o n   ( . % s )  U n s u p p o r t e d   c l i p b o a r d   f o r m a t  O u t   o f   s y s t e m   r e s o u r c e s  C a n v a s   d o e s   n o t   a l l o w   d r a w i n g # T e x t   f o r m a t   f l a g   ' % s '   n o t   s u p p o r t e d   ��ߘ{<:y&q?	*%TPF0TAboutDialogAboutDialogLeftuTop{HelpType	htKeywordHelpKeywordui_aboutBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	Om WinSCPClientHeight�ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenter
DesignSize�� PixelsPerInch`
TextHeight TButtonOKButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionOKDefault	ModalResultTabOrder OnMouseDownOKButtonMouseDown  TButtonLicenseButtonLeft>Top�WidthKHeightAnchorsakLeftakBottom Caption
&Licens...TabOrderOnClickLicenseButtonClick  TButton
HelpButtonLeftETop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelPanelLeft Top Width�Height�AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder
DesignSize��  TLabelApplicationLabelLeft>TopWidth4HeightCaptionApplicationShowAccelChar  TLabelVersionLabelLeft>TopWidthHeightCaptionVersion 2.0.0 (Build 12) XXShowAccelChar  TLabelWinSCPCopyrightLabelLeft>Top8Width� HeightCaption%   Copyright © 2000-2003 Martin PrikrylShowAccelChar  TLabelProductSpecificMessageLabelLeft>TopdWidthHeightCaption5   För att skicka in kommentarer och rapportera buggar:ShowAccelChar  TLabelLabel3Left>TopWidth[HeightCaption   Copyright för vissa delar:ShowAccelChar  TLabelRegistrationLabelLeft>Top� WidthHeightCaptionThis product is licensed to:ShowAccelChar  	TPaintBoxIconPaintBoxLeftTopWidth0Height0OnPaintIconPaintBoxPaint  TStaticTextHomepageLabelLeft>TopHWidth� HeightCaptionhttp://XXXXXXwinscp.net/TabOrder TabStop	  TStaticTextForumUrlLabelLeft>ToptWidth� HeightCaptionhttp://XXXXwinscp.net/forum/TabOrderTabStop	  TPanelThirdPartyPanelLeft>TopWidthRHeight� AnchorsakLeftakTopakRight 	BevelKindbkTile
BevelOuterbvNoneParentColor	TabOrder  TPanelRegistrationBoxLeft>Top� WidthRHeightYAnchorsakLeftakTopakRight 	BevelKindbkTile
BevelOuterbvNoneParentBackgroundParentColor	TabOrder
DesignSizeNU  TLabelRegistrationSubjectLabelLeftTopWidth� HeightAAnchorsakLeftakTopakRight AutoSizeCaptionSomeone
Somewhere, some cityShowAccelCharWordWrap	  TLabelRegistrationLicensesLabelLeftTop+WidthjHeightCaptionNumber of Licenses: XShowAccelChar  TStaticTextRegistrationProductIdLabelLeftTopAWidth� HeightCaptionProduct ID: xxxx-xxxx-xxxxxShowAccelCharTabOrder OnClickRegistrationProductIdLabelClick        TPF0TAuthenticateFormAuthenticateFormLeft0TopqHelpType	htKeywordHelpKeywordui_authenticateBorderIconsbiSystemMenu BorderStylebsDialogCaptionAuthenticateFormClientHeight|ClientWidthwColor	clBtnFaceConstraints.MinHeight� Constraints.MinWidth
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnResize
FormResizeOnShowFormShowPixelsPerInch`
TextHeight TPanelTopPanelLeft Top WidthwHeightAAlignalClient
BevelOuterbvNoneTabOrder  TListBoxLogViewLeft0Top WidthGHeightAStylelbOwnerDrawVariableAlignalClient
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneDoubleBuffered	ParentDoubleBufferedParentShowHintShowHint	TabOrder 
OnDrawItemLogViewDrawItemOnMeasureItemLogViewMeasureItemOnMouseMoveLogViewMouseMove  TPanel	LeftPanelLeft Top Width0HeightAAlignalLeft
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder 	TPaintBoxAnimationPaintBoxLeftTopWidth Height     TPanelPasswordPanelLeft TopAWidthwHeight� AlignalBottomAutoSize	
BevelOuterbvNoneTabOrderVisible TPanelPromptEditPanelLeft Top WidthwHeight� AlignalTop
BevelOuterbvNoneTabOrder 
DesignSizew�   TLabelInstructionsLabelLeftTopWidthhHeight'AnchorsakLeftakTopakRight AutoSizeCaption�Instructions for authentication. Please fill in your credentials carefully. Enter all required information, including your session username and session password.XFocusControlPromptEdit1WordWrap	  TLabelPromptLabel1LeftTop8WidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption&UsernameX:FocusControlPromptEdit1WordWrap	  TLabelPromptLabel2LeftTopeWidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption&PasswordX:FocusControlPromptEdit2WordWrap	  TPasswordEditPromptEdit1LeftTopIWidthiHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPasswordEditPromptEdit2LeftTopvWidthiHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPanelSavePasswordPanelLeft Top� WidthwHeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSavePasswordCheckLeftTopWidthHeightCaption   &Ändra lösenord till det härChecked	State	cbCheckedTabOrder    TPanelButtonsPanelLeft Top� WidthwHeight,AlignalTop
BevelOuterbvNoneTabOrder
DesignSizew,  TButtonPasswordOKButtonLeftvTopWidthKHeightAnchorsakTopakRight CaptionOKModalResultTabOrder   TButtonPasswordCancelButtonLeft� TopWidthKHeightAnchorsakTopakRight CaptionAvbrytModalResultTabOrder  TButtonPasswordHelpButtonLeft&TopWidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick   TPanelSessionRememberPasswordPanelLeft Top� WidthwHeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSessionRememberPasswordCheckLeftTopWidthHeightCaption.   &Kom ihåg lösenordet för den här sessionenChecked	State	cbCheckedTabOrder     TPanelBannerPanelLeft Top*WidthwHeightRAlignalBottom
BevelOuterbvNoneTabOrderVisible
DesignSizewR  TMemo
BannerMemoLeftTopWidthhHeight"AnchorsakLeftakTopakRightakBottom Color	clBtnFace	PopupMenuBannerPopupMenuReadOnly	
ScrollBars
ssVerticalTabOrder WantReturnsOnContextPopupBannerMemoContextPopup  	TCheckBoxNeverShowAgainCheckLeftTop5Width� HeightAnchorsakLeftakRightakBottom Caption&   &Visa aldrig det här meddelandet igenTabOrder  TButtonBannerCloseButtonLeft� Top/WidthKHeightAnchorsakRightakBottom Caption	   FortsättModalResultTabOrder  TButtonBannerHelpButtonLeft$Top/WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TActionList
ActionListLeft Top0 	TEditCopyEditCopyActionCategoryBannerCaptionK&opiera
ImageIndex ShortCutC@  TEditSelectAllEditSelectAllActionCategoryBannerCaption&Markera allt
ImageIndexShortCutA@  TActionBannerMonospacedFontActionCategoryBannerCaption   Använd typsnitt &Monospaced	OnExecute!BannerMonospacedFontActionExecute  TActionLabelCopyActionCategoryLabelCaptionK&opiera	OnExecuteLabelCopyActionExecute  TActionLabelOpenLinkActionCategoryLabelCaption   &Öppna	OnExecuteLabelOpenLinkActionExecute   
TPopupMenuBannerPopupMenuLeft� Top0 	TMenuItemCopyItemActionEditCopyAction  	TMenuItemSelectAllItemActionEditSelectAllAction  	TMenuItemN1Caption-  	TMenuItemAdjustWindowItemActionBannerMonospacedFontAction   
TPopupMenuLabelPopupMenuLeft8TopH 	TMenuItemCopy1ActionLabelCopyAction  	TMenuItemN2Caption-  	TMenuItemOpen1ActionLabelOpenLinkActionDefault	     TPF0TCleanupDialogCleanupDialogLeftdTop� HelpType	htKeywordHelpKeyword
ui_cleanupBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRensa applikationsdataClientHeight+ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize�+ PixelsPerInch`
TextHeight TLabelLabel1LeftTopWidth�HeightaAnchorsakLeftakTopakRight AutoSizeCaption8  Följande lista innehåller all data som det här programmet lagrar på den här datorn. Välj det som du vill ska tas bort.

Om ytterligare instanser av programmet är igång, var god avsluta dem innan nedanstående data tas bort.

Notera att en del av dessa data kommer att återskapas vid nästa uppstart.ShowAccelCharWordWrap	  TButtonOKButtonLeft� TopWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftITopWidthKHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  	TListViewDataListViewLeftTophWidth�Height� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsCaptionDataWidth�  CaptionPlatsWidth�  ColumnClickDoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowHint	TabOrder 	ViewStylevsReport	OnInfoTipDataListViewInfoTipOnKeyUpDataListViewKeyUpOnMouseDownDataListViewMouseDown  TButtonCheckAllButtonLeftTop
WidthqHeightAnchorsakLeftakBottom CaptionMarkera &allaTabOrderOnClickCheckAllButtonClick  TButton
HelpButtonLeft�TopWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick      TPF0TConsoleDialogConsoleDialogLeft]Top� HelpType	htKeywordHelpKeyword
ui_consoleBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionKonsolClientHeight�ClientWidth'Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth�
ParentFont		Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ' �'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�&!�                        '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�                        '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�                        '!�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�'!�                        '!�*$�*$�*$�*$�������������E@;�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�'!�                        '!�,% �,% �,% �2,'���������������������-&!�,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �'!�                        '!�.'!�.'!�.'!�.'!�������������������������TNI�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�'!�                        '!�0("�0("�0("�0("�;4.�����������������������������6.)�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�0("�'!�                        '!�2*$�2*$�2*$�2*$�2*$�2*$�c]X�������������������������f`\�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�2*$�'!�                        '!�4+%�4+%�4+%�4+%�4+%�4+%�4+%�80*�����������������������������@82�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�4+%�'!�                        '!�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�XQK�������������������������upk�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�'!�                        '!�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�80)�����������������������������JB<�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�7/(�'!�                        '!�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�OGA�������������������������~xt�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�'!�                        '!�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*��{v���������������������UMF�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�;2*�'!�                        '!�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+��zu���������������������WNG�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�'!�                        '!�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�ULE��������������������������{v�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�?5-�'!�                        '!�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�A7/�������������������������ÿ��TKD�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�'!�                        '!�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�bZS��������������������������ys�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�B8/�'!�                        '!�D91�D91�D91�D91�D91�D91�D91�H=6�����������������������������PE>�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�'!�                        '!�F;2�F;2�F;2�F;2�F;2�F;2�pga�������������������������umf�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�'!�                        '!�H<3�H<3�H<3�H<3�RF>�����������������������������NB9�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�'!�                        '!�J>5�J>5�J>5�J>5�������������������������lb[�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�'!�                        '!�K?6�K?6�K?6�PE<���������������������NB9�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�'!�                        '!�MA7�MA7�MA7�MA7�������������dYQ�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�MA7�'!�                        '!�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�'!�                        '!�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�'!�                        '!�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�'!�                        '!�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�UG<�'!�                        '!�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�VH>�'!�                        '!�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�'!�                        '!�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�'!�                        '!�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�\MB�'!�                        '!�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�'!�                        '!�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�'!�                        '!�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�aQF�'!�                        '!�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�'!�                        '!�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�eTH�'!�                        '!�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�'!�                        '!�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�iXK�'!�                        '!�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�'!�                        '!�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�l[M�'!�                        '!�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�n\O�'!�                        '!�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�'!�                        '!�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�'!�                        �] ��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��e'��] �                        �] ��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��w5��] �                        �] ��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��C��] �                        �] ��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��j��] �                        �] ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������] �                        �]ů] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��]�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ���������������������������������������������������������      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      ��������������������������������������������������������(   0   `          �%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�                '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�                '!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�'!�                '!�*$�*$�*$�������������/)#�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�*$�'!�                '!�-& �-& �-& �����������������]WS�-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �-& �'!�                '!�/("�/("�/("�tpl���������������������:4.�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�/("�'!�                '!�1*#�1*#�1*#�1*#�C<6���������������������qlg�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�'!�                '!�4,%�4,%�4,%�4,%�4,%�4,%�smh���������������������D<6�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�'!�                '!�6.'�6.'�6.'�6.'�6.'�6.'�6.'�A93����������������������|w�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�'!�                '!�90)�90)�90)�90)�90)�90)�90)�90)�90)�f_Z���������������������RKD�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�'!�                '!�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�@70���������������������=3,�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�'!�                '!�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�B81���������������������?5-�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�>4,�'!�                '!�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�kd]���������������������YPI�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�'!�                '!�C80�C80�C80�C80�C80�C80�C80�MC;�����������������������}�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�'!�                '!�E:2�E:2�E:2�E:2�E:2�E:2�wq���������������������UKC�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�E:2�'!�                '!�H<3�H<3�H<3�H<3�XMD�¾�������������������xr�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�H<3�'!�                '!�J>5�J>5�J>5��}w���������������������TH@�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�J>5�'!�                '!�M@7�M@7�M@7�����������������ukd�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�'!�                '!�OB9�OB9�OB9�������������SF=�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�OB9�'!�                '!�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�RD:�'!�                '!�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�'!�                '!�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�'!�                '!�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�YK@�'!�                '!�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�'!�                '!�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�^NC�'!�                '!�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�'!�                '!�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�'!�                '!�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�eUH�'!�                '!�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�'!�                '!�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�jYL�'!�                '!�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�m[N�'!�                '!�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�'!�                '!�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�'!�                �] ��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��] �                �] ��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��] �                �] ��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��Y��] �                �] ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������] �                �]��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��]�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������  ������  ������  ������  ������  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      ������  ������  ������  ������  ������  (   (   P          @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�        '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�        '!�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�("�'!�        '!�+$�+$�+$���������^XT�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�+$�'!�        '!�.'!�.'!�.'!�����������������93-�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�.'!�'!�        '!�1)#�1)#�1)#�6.(�����������������qkg�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�'!�        '!�4,%�4,%�4,%�4,%�4,%�WPJ�����������������G@9�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�4,%�'!�        '!�7.'�7.'�7.'�7.'�7.'�7.'�8/(������������������}y�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�7.'�'!�        '!�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�PHA�����������������:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�:1)�'!�        '!�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�SJC�����������������=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�=3+�'!�        '!�@6.�@6.�@6.�@6.�@6.�@6.�A7/�������������������|�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�@6.�'!�        '!�C80�C80�C80�C80�C80�cZT�������������¾��SIB�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�C80�'!�        '!�F:2�F:2�F:2�J>7�����������������wq�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�F:2�'!�        '!�I=4�I=4�I=4�����������������SG?�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�'!�        '!�K?6�K?6�K?6���������vmf�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�'!�        '!�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�NB8�'!�        '!�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�'!�        '!�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�TG<�'!�        '!�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�WI>�'!�        '!�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�'!�        '!�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�]NB�'!�        '!�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�'!�        '!�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�cSG�'!�        '!�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�'!�        '!�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�iWK�'!�        '!�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�lZM�'!�        '!�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�o\O�'!�        '!�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�r_Q�'!�        �] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] �        �] ��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��g)��] �        �] ��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��};��] �        �]��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��]�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �����   �����   �����   �����   �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �����   �����   �����   �����   (       @          �                                                                                                                                                                                                                                                                                      !!!!!!!!!!!!!!!!!!!!!!!!!!!!        '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�        '!�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�*#�'!�        '!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�.&!�'!�        '!�1*#�1*#�d^Y�����70*�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�1*#�'!�        '!�5-&�5-&�������������e_Z�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�5-&�'!�        '!�90)�90)�aZT�����������������D;4�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�90)�'!�        '!�=3,�=3,�=3,�A81�����������������{to�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�'!�        '!�A6.�A6.�A6.�A6.�A6.�bYR�����������������A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�'!�        '!�E:1�E:1�E:1�E:1�E:1�E:1���~�������������E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�E:1�'!�        '!�I=4�I=4�I=4�I=4�`VN�����������������`VN�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�I=4�'!�        '!�M@7�M@7�NA8���������������������M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�M@7�'!�        '!�PC9�PC9�������������¾��^RH�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�PC9�'!�        '!�TF<�TF<����������~w�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�TF<�'!�        '!�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�XJ?�'!�        '!�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�\MA�'!�        '!�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�`PD�'!�        '!�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�dSG�'!�        '!�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�gVJ�'!�        '!�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�kZL�'!�        '!�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�'!�        H*�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�uR8�H*�        p6��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0��p0�p6�        p6���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@�p6�        p6��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c��c�p6�        p6�����������������������������������������������������������������������������������������������������������������p6�        p5�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p5�                                                                                                                                                                                                                                                                                                                                                                                                    ���������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ������������(      0          `	                                                                                                                                                                                                                  ' �'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�,% �,% ���������/(#�,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �,% �'!�'!�1)#�1)#�KD?���������YSN�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�1)#�'!�'!�6.'�6.'�6.'�6.'���������>6/�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�6.'�'!�'!�<2+�<2+�ULF���������aXS�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�<2+�'!�'!�A6.�A6.���������B7/�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�A6.�'!�'!�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�F;2�'!�'!�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�'!�'!�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�QD:�'!�'!�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�VH=�'!�'!�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�[LA�'!�'!�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�'!�'!�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�fUI�'!�'!�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�kYL�'!�'!�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�p^P�'!��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��] ��] ��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��w��] ��] �] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] �                                                                                                                                                                                                ��� ���                                                                                 ��� ��� (      (          �                                                                                                                                                                                  '!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!���������.)$�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�'!�(!�ZTO���������\UQ�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�'!�'!�/'"�/'"�5-(�������������/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�'!�'!�6-'�6-'�90*�������������6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�'!�'!�=3,�bYS���������umg�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�'!�'!�D91���������ND<�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�D91�'!�'!�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�'!�'!�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�'!�'!�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�'!�'!�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�'!�'!�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�'!�'!�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�'!��] ��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��] ��] ��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��] ��] د] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] �                                                                                ��� ���                                                                     ��� (                 @                                                                                  '!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�' �'!�/'"�0(#�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�'!�'!�QIC�����slg�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�'!�'!�=3,�bYS���������QGA�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�'!�'!�D91�D91�RH@���������D91�D91�D91�D91�D91�D91�D91�D91�D91�'!�'!�L?6��vo���������SG>�L?6�L?6�L?6�L?6�L?6�L?6�L?6�L?6�L?6�'!�'!�i\S�����ui`�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�'!�'!�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�'!�'!�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�'!�'!�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�'!�'!�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�'!��] ��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��s2��] ��] ��w��w��w��w��w��w��w��w��w��w��w��w��w��w��] ��] د] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] ��] �                                                                ��                                                          ��  OldCreateOrder	OnCloseQueryFormCloseQueryOnShowFormShow
DesignSize'� PixelsPerInch`
TextHeight TBevelBevel1Left Top Width'HeightNAlignalTopShapebsBottomLine  TLabelLabel1Left3TopWidthNHeightCaptionAnge &kommando:FocusControlCommandEdit  TLabelLabel2Left3Top8WidthWHeightCaptionAktuell katalog:ShowAccelChar  TLabelLabel4Left3Top"Width�HeightAnchorsakLeftakTopakRight AutoSizeCaptionP   Varning: Kör inga kommandon som kräver användardata eller dataöverföringar.ShowAccelChar  
TPathLabelDirectoryLabelLeft� Top8Width+HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TImageImageLeftTopWidth Height AutoSize	  TMemo
OutputMemoLeft TopNWidth'Height;TabStopAlignalClientColor	clBtnFace	PopupMenu	PopupMenuReadOnly	
ScrollBarsssBothTabOrderWantReturnsOnContextPopupOutputMemoContextPopup  TButton	CancelBtnLeft�TopWidthKHeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  THistoryComboBoxCommandEditLeft� Top	Width� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength TabOrder OnChangeCommandEditChange  TButtonExecuteButtonLeft�TopWidthKHeightAnchorsakTopakRight Caption   K&örDefault	TabOrderOnClickExecuteButtonClick  TButton
HelpButtonLeft�Top*WidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPngImageListImages	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?Cf���X�1&���Ӳþ`��e=��(�g���?���K��t���VC��w��?�,����(
>}��p��+���/�a`f�U����k�Ϫf(�u .�o��������W�+�_1��u�����������_�D��m؃-L�$���?�*��t�A����>2`�#�2�ه�I�+�Ϫg��₪i���Ʌs̬�3�}ހHhZ�vu$C�\�>��0�<g�\����Wg���oX�vMû���k�md@8���kO��;�1 �l@\����j���K~x��9LЁ��æ�g�V�A��]4 ������c@t�����i��F@������Y�����GZ3���fXP1���EA\��0�jH�*������]�&�(̊��o%â�X�D�,@	l��9Ò�x�DU���@Xښ� Ld8��h��    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�d@D�l�LYљ�7`ak
I�����%C���������́!�P3Հy�.�z°x�1�7�?��|<�����z�p5I�h�mJ����7Cq�
���2ؙh0�����ȹ[l�,��bX������0�b��_�n�����Ƞ�&����?���k�~���W�Nj=��������ÉKwn���%��o?��]��\`vZ�3�!|����y��o� �W�c�T�b�y���%d4�0�.,q��u�U�O0��3D�X�Ū&�b���+Cgq$܀����L��p��=��2�
�1��2\�������`���`1a>0;�̀�5	`���x��b7��  +!� "��p���hkU�xn�T&A �(��������e���8*��X�j���X�0��ߊf E��  O	��NV    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  2IDATx�c���?�y�u��mF���JI�=���n��M��:�b����O���/�g�+�*w��v���N
�,�g�Dfa�_<�a�����εs04����?�0@M�,�w�bg�X�"|�[WN#PT�c8�cX��#�$�·�����n`8��9 �>�w�<P� 	iE�Ӈ��%Lm1C��Լxza���4X���p��o_=E�'(�⼫g�`8Y�5�>��0���C��˧�lu]S�o_?#`ecg��ݸȠ���U����p>�<��/`( �h����`    IEND�B`�  LeftHTop� Bitmap
      
TPopupMenu	PopupMenuImagesImagesLeft�Top�  	TMenuItemCopyItemActionEditCopy  	TMenuItemSelectAllItemActionEditSelectAll  	TMenuItemN1Caption-  	TMenuItemAdjustWindowItemActionAdjustWindow   TActionList
ActionListImagesImages	OnExecuteActionListExecuteOnUpdateActionListUpdateLeftHTop�  	TEditCopyEditCopyCaptionK&opiera
ImageIndex ShortCutC@  TEditSelectAllEditSelectAllCaption&Markera allt
ImageIndexShortCutA@  TActionAdjustWindowCaption   Anpassa &fönster
ImageIndexShortCutJ@   TPngImageList	Images120HeightWidth	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  CIDATxڍ��ORaǿgm���П�}��m��&3�����]t�px�rfkp	���R��njβ�[s���EƜ�&F
�	��Ǿgg;�����|vG��#���*�	QWd��Y�����i�q
�mB����*s�7�R��^�3E�,(��P��e|\]�����(��%��1�'�d���bא�t��!�/)����rȦ�0��IH�D����0���§o��Jza�i�	<�?ABvn��,�d5�fo��N=�mՂ#�,Ys�Ҙ��Д��xbu ��nX���^�R�,�Ko�r��P�!� M�(�]<6�����GV�]����~@�.ᗪ�͍X�>G�K�)K:9��&��녚jA<MVk�k���"�]htܫ74��W��d��T���Fĥo y!BBb2[Uՠ70	���XGa�'u���&I4#���
<M���hl ���o��� h�ZsMw�o�=g@��~I0:�TY��1�xMl o�Pe���0�F�ϱ�[�*��/�؀��y�4Y���#�����HdO�?�^���f���� m    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  CIDATx�c���?5#�����T1uEg*#����)_=��-��P3���h~���aݞ��n=ax��XL���AWU�!�̈́���E}"��������m�f�G��bu��� CSv 33\,����M����x�Q0[_]���P���.0��qmE����8\Or��s����^�c�~�óWb},XX����O]gX��8����`��דR?��YH"���1<}�����'/ޅCr�=���2\]��3P�q�9Þ�Wn ]���_���PLo@3pF=��S��2�[w�fzWCQ�A]Q����_[]�x1ؑ����hN�O�K6O� ��`�곃�x�����fX����(f6�G5pZ���� q~^.���pFF����N_�Iw@/��(��d5�8�a`��u/�|����Ud.�|�p����/+[cu$G�8���W�1,\#"�5�.�xf��0�����r��\����������DyLu���<r����_l���p��-P�X��@	�oE3pBe��H�iP 7��  J�I�^�D+    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
`  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?5�B��@Z�J���?�׉*��ܼ���Bb2x�;J���_�U���FE���68y;3ą��ًVnfX�u/N�g���g�UA��CbT ���e��lڅU��S�!jX��ʮu���[P^u�/���e��aX�v���[��iG�h9d=w���(�������`����Ȯ5`���9K������������9�8�b���O؂S͔��:;;!�471�G��Tld�
��ۍS�¥�jj� 
�1�e0$�E1��a(�|���%7o�2��I3>�{1���,YR����?CӍK'����9����_>Bdc�`��޸ ��5�����@`�UAUy	Cfz2����s�:{p�f n 14j�<�A Aa�� !��J+�z���J" �e_�^bS�@ ����;e*    IEND�B`�  Left�Top� Bitmap
      TPngImageList	Images144HeightWidth	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  rIDATxڵ��KSaƯ}�/I����0�,�(�R�e-��5�4�*綳��NLTf�IBQ��K	"(���M�mns�ŧg��v�?x}<���;7��B��EWL�X(oa�e9^��hwpW��c�����w�~��$�� �?dj΁��U�~�1A�L�r��Ն��^�>B��k�A�λ�����}����,f��{AԲ\����J���n����KD0�}��D̀*�i�ʇ7\ؠ�˞5�-����ZlD+/���8�}ŗ�/�LK *�]u\�pڭ_n/��Sجi	���Jt5G�Y'�.��X��d�3j��m?d�f/� �,��=�eZ�.+nڟ@&��� �\TgOT�i:����!\}1���,��جi��\QpZ��试bq���f��MsS�������j� �B�v�{��9W�ɴ?);�
���� ��6�]?�'�.zA�S꾀i�i0�PS��=��r8W����2-9�]P�Sݱ��LK۶i�Qr�hS��D��_=ʚ�MK�q�T�0+�� ��SдԨ�t6I��
��i�9�w'5��Y�(�H������=�+�ŵ&A�RӤ�Bo������� le~���v�h    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
/  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-#�,�(�M5�Vt�2b�`ak
ņ�W��m���d�-H���ۂ�h������p����o>2|�񋁃��AB����@���B���ՂD|�kF�`ƪ��.���ZkCU�� ;��Z<�mBXp����E;�lf&S]%N�{O^1�}�
���$�A���O��c���$����2<}�������f��`+�[����0�$ѓACQ�/�nnf7",@��&&��w�2LZ�����`~v����\}j=f5`Z���7pp�~���0h^���"���`����7�`&����gX������pq6V�o~����Ǻ3h)K����Y0�>�p��[��y�8�L��)J�2LZ������b�4����2��`z�I��~�DdQ�'���\�{�Vpp�@�%��Mx,��dAN�BxД��2�K�@#�C��u�����8AOM�/�Sk�������;0[\����F������}��ӗ�pu�~��*p~v3&�$�^��a�������AMA��ƽ�`���6C��)\>�en&!Y �n>b�u���o��GUA�}p���v�����!���'��(��x,�PE�mx,��t(�j��з  �n���    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  `IDATx�c���?-#�-P�]� H����� ���:�������}�_HL�&�{�b��e��������QFQ����'A�Ғb}M%`vQ]����9sx;��
���&��3�H���O��d(��d���^}N�X�kb�WaIN"����ؾC'z��ǫ��4��
�]��i��$��_�pb���	"8��
�:�gbhطy	�v���+/Lg�0m>�ϟ�`�}��Eu}����4CKm1����0����`����Oj�{�4ܿyb������#Ci^:����k�>�{N5 tO�ɰ}�~�Gw�A,��Sa��pz3h;N��>`��-x,�	�i[w�ex���1)HQ�(/���V�e�m�14�=�L㒻��1CiU�~{��!�!Q)�Bv���ڦNC.�����1ˮ�r�֮	?~����{�b��(1����`Z�ؖ(�߿�X��ˏWagk��jq�q�v������~������B�Mk�1()*����?`�����~��������w���lXf��1ܽw���?~C, *@� 8�L�]��X-@ԟ202H��4����>�-  �+�`{O�    IEND�B`�  LeftHTop Bitmap
      TPngImageList	Images192Height Width 	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�ŕ�OQ�O7�����q�QB���>���n4
h��C5B�
��"��QQ	$�� 5<
�o�-ס!���tF��������L�W	!��6��G��$!�d5���J�����w Jt/I��3�S��#�C��:7o05Y*����r�,"�����'�ѩ�c˾PjoT��/���9�G�|�sa��k5���_H �f�*\����'���7`x>�:���1x�!,��� �x?13m*��"�j�3�@�O�WS�1�y����>�
���� �NbVe�����D��{��a�}!���Ck�%� W��\!�'�u�v6��3��0;��Z�) ��N,U2���>�(N?[��h�ȅ��� V�W<~4�}J�!��� 9�.bQ+��gp�PG�#xע+,*@��)�h���O܀�Os�(�
�
���` �����>La��=
��2V�]q ��6b������o ��
�ٟ�PY�I���:�]�ԁ�hA���
�ٿs[v ��b��a����U���-�
ˢʈ�����:�Lf������+��J)@�a�7`vA���j�I�����g\�bK����1�� 0t����HO��2�Z%�Ϡ�KXlQ5��I��x �����U�¢�Dvr@׍��� �
+���R����.O8����SX�+O�Vu���|� ��.a�E��D��� ��&Na�R(;[����P ���r�� �֞p	k���+T���_6��/�.    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  rIDATx���{PLQ�o�^[D�d*=��#�h��c�ь�fL驄J�0���˫H��P�͘A�`H�I[
���d%=��������=�=�?~�����9�{ν�h����_���"�g�ٿ��9�1&�bb�Z'��9����V�֘�܀����� 29 �}b���m+�;����Y����0�l;�iX��^�+��C�5B�^)@�x��	y���񀽍�j�
 C@�كؔ[��2��h#9���i��	$ �j*���&�ϱ���!��Q��
�����:7���c�R �Y%�L�����ɅnZ+�-��W�����-Y8~�n 86�p�` �iH:ys{'�?���+֯X@�d�)���:����!��D]H�o �B��u�6�VB�*b���e���}�P�؆���h� h��g4��LG��j"�-�83�U��
��FzSWfޜۼ�ȇ� iq$���	��
�˭�<�Y��KO�B&����܉���T@ ���3�{4W�;S&����=�f[��P_���_����J��* �܀�J���d�~̴x����}��.�n)��Ǵ" H`;p*��v�Ee�L����[��tO�m,@�	O� R� 7��QXZôyz:H�����ӂ���PK�=��=�*� �F���Ŭ���1V�9A[k�_7�Ie=�eؘ� �-	8D�(�$ĝ��.�[�:�Z��Jv%��!�v� '����'\��|֗�榓�q���X5{C<1�ĈU��p7��
�,dw@�ӗ�{'��^�;0m�D,r����LhH�|PR�
������]P�* F5�OED"p\̀H��>���( ���#��������H��    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�c���?�@�Q����#�*]m��p��� 5��6�ϊt���Ӗ�a��(�� �:�Ε������|z�p����S[/�q�6���!Y����߻�p���I�H�3����م5]O��$I��c�P�o�D�fv66���`G� ����v���~m�œ�P�kbO�撜D';�D���	��)�6�򙃨�2�&)A`�ڹ`�=8�d���Eu���9Ɇ�ٰL�ē��楓�P�6!ِ}���i'���޾z�JpIvv6������ix9�m��������(��o���?��ލ��W�K���0�Օ2��J3ظ��5���5`�u?e�j�fx��	X���+��U�`�rsb(-� � 1��9 Lۻ�(���0�a�.`��Rr*���Y@�e����>y`�����?�a뎽��Au���"X���,Cwk-��6���k�����41�<|�PZ��pH��˧�Q *!�����PY��P�҅��s�v�i#+W��k��{&2���.���cT�J������`Z�ܑd��^?Gu ��(Ɇ\9sL�ؒ���ר��'�=p��10�ihE��/ߡ:����h�]m��>�	o��eU�D����'T�sp�����a��eJ�
`����������f��������}PVRdؼR�F0ܽw�$���Du 3I�@P��^�a�z����� �M�@8@Q�#�2]m������7UG�lD;  �/���J{�    IEND�B`�  Left�Top Bitmap
       TPF0TCopyDialog
CopyDialogLeftkTop� HelpType	htKeywordHelpKeywordui_copyBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
CopyDialogClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight TImageImageLeftTopWidth Height AutoSize	  TLabelDirectoryLabelLeft.TopWidth� HeightCaption)Copy 2 selected files to remote directory  THistoryComboBoxLocalDirectoryEditLeft.TopWidthtHeightAutoCompleteAnchorsakLeftakTopakRight DropDownCountTabOrder TextLocalDirectoryEditOnChangeControlChangeOnExitLocalDirectoryEditExit  THistoryComboBoxRemoteDirectoryEditLeft.TopWidth�HeightAutoCompleteAnchorsakLeftakTopakRight DropDownCount	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  TButtonOkButtonLeftTop� WidthKHeightAnchorsakTopakRight CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftWTop� WidthKHeightAnchorsakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonLocalDirectoryBrowseButtonLeft�TopWidthKHeightCaption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick  	TCheckBoxQueueCheck2LeftToppWidth=HeightCaption1Transfer on background (add to transfer &queue) XTabOrderOnClickControlChange  TButton
HelpButtonLeft�Top� WidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  	TCheckBoxNeverShowAgainCheckLeftTop� Width�HeightCaption$   &Visa inte den här dialogrutan igenTabOrder
OnClickNeverShowAgainCheckClick  TButtonTransferSettingsButtonLeftTop� Width� HeightCaption   Överförin&gsinställningar...StylebsSplitButtonTabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxCopyParamGroupLeftTop5Width�Height2Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamGroupClick   TPanelShortCutHintPanelLeft Top� Width�Height"AlignalBottom
BevelOuterbvNoneParentBackgroundTabOrder	 TLabelShortCutHintLabelLeftTopWidth�HeightAutoSizeCaption�   I Commander-gränssnittet används kortkommandot F5 för att överföra filer. Om du vill använda kommandot för att uppdatera en filpanel, klicka här för att gå till inställningar.ShowAccelCharWordWrap	OnClickShortCutHintLabelClick       TPF0TCopyParamCustomDialogCopyParamCustomDialogLeftvTop� HelpType	htKeywordHelpKeywordui_transfer_customBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption   ÖverföringsinställningarClientHeightClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQuery
DesignSize� PixelsPerInch`
TextHeight TButtonOkButtonLeft� Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  �TCopyParamsFrameCopyParamsFrameLeft Top Width�Height�HelpType	htKeywordTabOrder   TButton
HelpButtonLeftPTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0TCopyParamPresetDialogCopyParamPresetDialogLeftTopzHelpType	htKeywordHelpKeywordui_transfer_presetBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCopyParamPresetDialogClientHeight0ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�0 PixelsPerInch`
TextHeight TLabelLabel1Left
TopWidthZHeightCaption   Förinställnings&beskrivningFocusControlDescriptionEdit  TButtonOkButtonLeft�TopWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft�TopWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TEditDescriptionEditLeft
TopWidth�Height	MaxLength� TabOrder OnChangeControlChange  �TCopyParamsFrameCopyParamsFrameLeftTop3Width�Height�HelpType	htKeywordTabOrder  	TGroupBox	RuleGroupLeft�Top[Width� Height�AnchorsakLeftakTopakRightakBottom Caption   Regler för automatiskt valTabOrder
DesignSize� �  TLabelLabel2LeftTopWidthOHeightCaption   Mask värdna&mnFocusControlHostNameEdit  TLabelLabel3LeftTopDWidthOHeightCaption   Mask an&vändarnamnFocusControlUserNameEdit  TLabelLabel4LeftToptWidthrHeightCaption   Mask &fjärrkatalogFocusControlRemoteDirectoryEdit  TLabelLabel5LeftTop� WidtheHeightCaptionMask &lokal katalogFocusControlLocalDirectoryEdit  TEditHostNameEditLeftTop$Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnExitMaskEditExit  TEditUserNameEditLeftTopTWidth� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditRemoteDirectoryEditLeftTop� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditLocalDirectoryEditLeftTop� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TButtonCurrentRuleButtonLeftTop� WidthIHeightCaptionAktuellTabOrderOnClickCurrentRuleButtonClick  TStaticTextRuleMaskHintTextLeft_Top� Width� Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionMasktipsTabOrderTabStop	   	TCheckBoxHasRuleCheckLeft�TopBWidth� HeightAnchorsakLeftakTopakRight Caption'   Välj automatiskt förinställning närTabOrderOnClickControlChange  TButton
HelpButtonLeftOTopWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TCopyParamsFrameCopyParamsFrameLeft Top Width�Height�HelpType	htKeywordTabOrder  	TGroupBoxCommonPropertiesGroupLeft� Top� Width� HeightyCaption
AlternativTabOrder
DesignSize� y  TLabelSpeedLabel3LeftTop]WidthBHeightCaption&Hastighet (kB/s)FocusControl
SpeedCombo  	TCheckBoxPreserveTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Behåll tidsstä&mpelParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxCommonCalculateSizeCheckLeftTopCWidth� HeightAnchorsakLeftakTopakRight Caption   B&eräkna total storlekParentShowHintShowHint	TabOrderOnClickControlChange  THistoryComboBox
SpeedComboLeftjTopZWidthUHeightAutoCompleteTabOrderText
SpeedComboOnExitSpeedComboExitItems.Strings	Unlimited10245122561286432168   	TCheckBoxPreserveTimeDirsCheckLeft Top,Width� HeightAnchorsakLeftakTopakRight CaptionInklusive katalogerParentShowHintShowHint	TabOrderOnClickControlChange   	TGroupBoxLocalPropertiesGroupLeft� TopWidth� Height2CaptionNedladdningsalternativTabOrder
DesignSize� 2  	TCheckBoxPreserveReadOnlyCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Behåll skrivsky&ddParentShowHintShowHint	TabOrder    	TGroupBoxRemotePropertiesGroupLeftTop� Width� Height� Caption   ÖverföringsalternativTabOrder 	TCheckBoxPreserveRightsCheckLeftTopWidth� HeightCaption   Sätt fil&rättigheterParentShowHintShowHint	TabOrder OnClickControlChange  
TComboEdit
RightsEditLeft"Top,Width{Height
ButtonHint   Konfigurera filrättigheterClickKey@ParentShowHintShowHint	TabOrderText
RightsEditOnButtonClickRightsEditButtonClickOnExitRightsEditExitOnContextPopupRightsEditContextPopup  	TCheckBoxIgnorePermErrorsCheckLeftTopIWidth� HeightCaption   Ign&orera filrättighetsfelParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxClearArchiveCheckLeftTop`Width� HeightCaptionRensa 'Arki&v' attributTabOrder  	TCheckBoxRemoveCtrlZAndBOMCheckLeftTopwWidth� HeightCaptionRemo&ve BOM and EOF marks XTabOrderOnClickControlChange  	TCheckBoxEncryptNewFilesCheckLeftTop� Width� HeightCaption&Kryptera nya filerTabOrderOnClickControlChange   	TGroupBoxChangeCaseGroupLeftTopWidth� Height� Caption   Ändra filnamnTabOrder
DesignSize� �   TRadioButtonCCLowerCaseShortButtonLeftTopZWidth}HeightAnchorsakLeftakTopakRight CaptionGemener &8.3TabOrder  TRadioButtonCCNoChangeButtonLeftTopWidth}HeightAnchorsakLeftakTopakRight Caption   I&ngen förändringTabOrder   TRadioButtonCCUpperCaseButtonLeftTop,Width}HeightAnchorsakLeftakTopakRight Caption	&VersalerTabOrder  TRadioButtonCCLowerCaseButtonLeftTopCWidth}HeightAnchorsakLeftakTopakRight Caption&GemenerTabOrder  	TCheckBoxReplaceInvalidCharsCheckLeftTopqWidth}HeightCaption   &Ersätt '\:*?' ...TabOrderOnClickControlChange   	TGroupBoxTransferModeGroupLeftTopWidth� Height� Caption   ÖverföringslägeTabOrder 
DesignSize� �   TLabelAsciiFileMaskLabelLeftTopZWidth� HeightAnchorsakLeftakTopakRight Caption'   Överför följande &filer i textläge:FocusControlAsciiFileMaskCombo  TRadioButtonTMTextButtonLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption&Text (text, html, skript, ...)TabOrder OnClickControlChange  TRadioButtonTMBinaryButtonLeftTop,Width� HeightAnchorsakLeftakTopakRight Caption   &Binärt (arkiv, doc, ...)TabOrderOnClickControlChange  TRadioButtonTMAutomaticButtonLeftTopCWidth� HeightAnchorsakLeftakTopakRight Caption&AutomatisktTabOrderOnClickControlChange  THistoryComboBoxAsciiFileMaskComboLeftTopjWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextAsciiFileMaskComboOnExitValidateMaskComboExit   	TGroupBox
OtherGroupLeftTopRWidth�Height� Caption   ÖvrigtTabOrder
DesignSize��   TLabelIncludeFileMaskLabelLeftTopWidth/HeightCaptionFilmas&kFocusControlIncludeFileMaskCombo  THistoryComboBoxIncludeFileMaskComboLeftTop$Width&HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextIncludeFileMaskComboOnExitValidateMaskComboExit  TButtonIncludeFileMaskButtonLeft;Top!WidthPHeightCaption&Redigera...TabOrderOnClickIncludeFileMaskButtonClick  	TCheckBoxNewerOnlyCheckLeftTopOWidth� HeightCaption!Endast &nya och uppdaterade filerParentShowHintShowHint	TabOrderOnClickControlChange  TStaticTextIncludeFileMaskHintTextLeft� Top:Width}Height	AlignmenttaRightJustifyAutoSizeCaptionmasktipsTabOrderTabStop	  	TCheckBoxExcludeHiddenFilesCheckLeft� TopOWidth� HeightCaptionExkludera &dolda filerParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxExcludeEmptyDirectoriesCheckLeftTopfWidth� HeightCaptionE&xkludera tomma katalogerParentShowHintShowHint	TabOrderOnClickControlChange      TPF0TCreateDirectoryDialogCreateDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeywordui_create_directoryBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSkapa katalogClientHeight� ClientWidthQColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizeQ�  PixelsPerInch`
TextHeight TLabel	EditLabelLeftTopWidthUHeightCaptionNytt &katalognamn:FocusControlDirectoryEdit  TEditDirectoryEditLeftTopWidthAHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextDirectoryEditOnChangeDirectoryEditChange  TPanel	MorePanelLeft Top2WidthQHeight� AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSizeQ�   	TGroupBoxAttributesGroupLeftTopWidthBHeight� AnchorsakLeftakTopakRightakBottom Caption
EgenskaperTabOrder  �TRightsFrameRightsFrameLeftTop$Width� HeightWTabOrder �	TCheckBoxDirectoriesXCheckVisible   	TCheckBoxSetRightsCheckLeftTopWidth� HeightCaption   Sätt fil&rättigheterParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTop� Width-HeightCaption*   Använd &samma inställningar nästa gångTabOrder    TButtonOKBtnLeft[Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0TCustomCommandDialogCustomCommandDialogLeft�Top� HelpType	htKeywordHelpKeywordui_customcommandBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCustomCommandDialogClientHeight5ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�5 PixelsPerInch`
TextHeight 	TGroupBoxGroupLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize�  TLabelDescriptionLabelLeftTopWidth9HeightAnchorsakLeftakTopakRight Caption&BeskrivningFocusControlDescriptionEdit  TLabelLabel1LeftTop@WidthXHeightAnchorsakLeftakTopakRight Caption&Eget kommando:FocusControlCommandEdit  TLabelShortCutLabelLeftTop� Width]HeightCaptionKor&tkommando:FocusControlShortCutCombo  TEditDescriptionEditLeftTop WidthzHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  THistoryComboBoxCommandEditLeftTopPWidthzHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength TabOrderOnChangeControlChange	OnGetDataCommandEditGetData	OnSetDataCommandEditSetData  	TCheckBoxApplyToDirectoriesCheckLeftTop� Width� HeightCaption   &Tillämpa på katalogerTabOrderOnClickControlChange  	TCheckBoxRecursiveCheckLeft� Top� Width� HeightCaption   Kör &rekursivtTabOrderOnClickControlChange  TRadioButtonLocalCommandButtonLeft� TopzWidth� HeightCaption&Lokalt kommandoTabOrderOnClickControlChange  TRadioButtonRemoteCommandButtonLeftTopzWidth� HeightCaption   &FjärrkommandoTabOrderOnClickControlChange  	TCheckBoxShowResultsCheckLeftTop� Width� HeightCaption!   &Visa resultat i terminalfönsterTabOrderOnClickControlChange  	TCheckBoxCopyResultsCheckLeftTop� Width� HeightCaption&Kopiera resultat till urklippTabOrder	OnClickControlChange  TStaticTextHintTextLeftTopgWidthuHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  	TComboBoxShortCutComboLeft� Top� Width� HeightTabOrder
  	TCheckBoxRemoteFilesCheckLeft� Top� Width� HeightCaption   &Använd fjärrfilerTabOrderOnClickControlChange   TButtonOkButtonLeft� TopWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� TopWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftLTopWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TCustomDialogCustomDialogLeft�Top� BorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSave session as siteXClientHeight)ClientWidthFColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenter
DesignSizeF) PixelsPerInch`
TextHeight TButtonOKButtonLeftDTop	WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top	WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder   TButton
HelpButtonLeft� Top	WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TCustomScpExplorerFormCustomScpExplorerFormLeft� Top� CaptionCustomScpExplorerFormClientHeight�ClientWidthlColor	clBtnFace
ParentFont	
KeyPreview	OldCreateOrderOnClose	FormCloseOnCloseQueryFormCloseQueryOnConstrainedResizeFormConstrainedResizeOnShowFormShowPixelsPerInch`
TextHeight 	TSplitterQueueSplitterLeft Top!WidthlHeightCursorcrSizeNSHintR   Dra för att ändra storlek på kölistan. Dubbelklicka för att dölja kölistan.AlignalBottomAutoSnapMinSizeFResizeStylersUpdateOnCanResizeQueueSplitterCanResize  TTBXDockTopDockLeft Top WidthlHeight	FixAlign	  TPanelRemotePanelLeft TopWidthlHeightAlignalClient
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder  	TSplitterRemotePanelSplitterLeft� Top Height� CursorcrSizeWEAutoSnapMinSizeFResizeStylersUpdate  TTBXStatusBarRemoteStatusBarLeft Top� WidthlHeightPanels ParentShowHintShowHint	UseSystemFontOnClickRemoteStatusBarClickOnMouseDownRemoteStatusBarMouseDown  TPanelRemoteDirPanelLeft� Top Width�Height� AlignalClient
BevelOuterbvNoneTabOrder TUnixDirViewRemoteDirViewLeft Top Width�Height� AlignalClientDoubleBuffered	FullDrag	HideSelectionParentDoubleBuffered	PopupMenu&NonVisualDataModule.RemoteDirViewPopupTabOrder 	ViewStylevsReportOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterRemoteDirViewEnterOnExitDirViewExit	OnKeyDownDirViewKeyDown
OnKeyPressDirViewKeyPressOnResizeRemoteDirViewResize
NortonLikenlOffUnixColProperties.ExtWidthUnixColProperties.TypeVisibleOnDDDragFileNameRemoteFileControlDDDragFileNameOnBusyDirViewBusyOnChangeFocusDirViewChangeFocusOnSelectItemDirViewSelectItemOnLoadedDirViewLoaded
OnExecFileDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDDragDetectRemoteFileControlDDDragDetectOnDDEndRemoteFileControlDDEndOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectOnContextPopupRemoteDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnDisplayPropertiesRemoteDirViewDisplayPropertiesOnReadRemoteDirViewRead  TTBXToolbarReconnectToolbarLeft� ToppWidthkHeightCaptionReconnectToolbarImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem254Action*NonVisualDataModule.ReconnectSessionAction    TPanelRemoteDrivePanelLeft Top Width� Height� AlignalLeft
BevelOuterbvNoneTabOrder TUnixDriveViewRemoteDriveViewLeft Top Width� Height� DirViewRemoteDirViewOnDDDragFileNameRemoteFileControlDDDragFileNameOnDDEndRemoteFileControlDDEndUseSystemContextMenuOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDDragDetectRemoteFileControlDDDragDetectOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectAlignalClientDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedReadOnly	TabOrder OnEnterRemoteDriveViewEnterOnBusyDirViewBusy    TPanel
QueuePanelLeft Top$WidthlHeight� AlignalBottom
BevelOuterbvNoneTabOrder 
TPathLabel
QueueLabelLeft Top WidthlHeightIndentVerticalAutoSizeVertical	OnGetStatusQueueLabelGetStatusAutoSizeTransparent  	TSplitterQueueFileListSplitterLeft TopuWidthlHeightCursorcrSizeNSHintd   Dra för att ändra storlek på köfilens lista. Dubbelklicka för att dölja listan över köfiler.AlignalBottomAutoSnapMinSize
ResizeStylersUpdateOnCanResizeQueueFileListSplitterCanResize  	TListView
QueueView3Left Top-WidthlHeightHAlignalClientColumnsCaption	OperationWidthF Caption   KällaWidth�  Caption   MålWidth�  	AlignmenttaRightJustifyCaption
   ÖverförtWidthP 	AlignmenttaRightJustifyCaptionTidWidthP 	AlignmenttaRightJustifyCaption	HastighetWidthP 	AlignmenttaCenterCaption
UtvecklingWidthP  ColumnClickDoubleBuffered	DragModedmAutomaticReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuNonVisualDataModule.QueuePopupSmallImagesGlyphsModule.QueueImagesStateImagesGlyphsModule.QueueImagesTabOrder 	ViewStylevsReportOnChangeQueueView3ChangeOnContextPopupQueueView3ContextPopup
OnDeletionQueueView3DeletionOnEnterQueueView3EnterOnExitQueueView3Exit
OnDragDropQueueView3DragDrop
OnDragOverQueueView3DragOverOnSelectItemQueueView3SelectItemOnStartDragQueueView3StartDrag  TTBXDock	QueueDockTagLeft TopWidthlHeight	AllowDrag TTBXToolbarQueueToolbarLeft Top CaptionQueueToolbarImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder  TTBXItemQueueEnableItemAction%NonVisualDataModule.QueueEnableAction  TTBXSeparatorItemTBXSeparatorItem203  TTBXItem
TBXItem201Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem
TBXItem202Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem
TBXItem203Action)NonVisualDataModule.QueueItemPromptAction  TTBXItem
TBXItem204Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem195Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem194Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem
TBXItem205Action)NonVisualDataModule.QueueItemDeleteAction  TTBXSeparatorItemTBXSeparatorItem201  TTBXItem
TBXItem206Action%NonVisualDataModule.QueueItemUpAction  TTBXItem
TBXItem207Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem57  TTBXItem"QueueDeleteAllDoneQueueToolbarItemAction,NonVisualDataModule.QueueDeleteAllDoneAction  TTBXSeparatorItemTBXSeparatorItem202  TTBXSubmenuItemTBXSubmenuItem27Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem211Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem225Action3NonVisualDataModule.QueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem173Action0NonVisualDataModule.QueueSuspendOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem226Action1NonVisualDataModule.QueueShutDownOnceEmptyAction2	RadioItem	   TTBXItem
TBXItem208Action*NonVisualDataModule.QueuePreferencesAction    	TListViewQueueFileListLeft TopxWidthlHeightAlignalBottomColumns  DoubleBuffered		OwnerData	ReadOnly	ParentDoubleBufferedShowColumnHeadersTabOrderTabStop	ViewStylevsReportOnCustomDrawItemQueueFileListCustomDrawItemOnDataQueueFileListDataOnEnterQueueFileListEnterExitOnExitQueueFileListEnterExitOnResizeQueueFileListResize   TThemePageControlSessionsPageControlLeft Top	WidthlHeight
ActivePage	TabSheet1AlignalTopDoubleBuffered	ParentDoubleBufferedTabOrderTabStopOnChangeSessionsPageControlChangeOnContextPopupSessionsPageControlContextPopup
OnDragDropSessionsPageControlDragDrop
OnDragOverSessionsPageControlDragOverOnMouseDownSessionsPageControlMouseDownOnCloseButtonClick#SessionsPageControlCloseButtonClick 	TTabSheet	TabSheet1Caption	TabSheet1   TApplicationEventsApplicationEventsOnDeactivateApplicationEventsDeactivate
OnMinimizeApplicationMinimizeOnModalBeginApplicationEventsModalBegin	OnRestoreApplicationRestoreLeftXTop�    TPF0TEditMaskDialogEditMaskDialogLeftqTopHelpType	htKeywordHelpKeywordui_editmaskBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRedigera filmaskClientHeight�ClientWidth�Color	clBtnFace
ParentFont	
KeyPreview	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBox
FilesGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption	FilmaskerTabOrder 
DesignSize��   TLabelLabel3LeftTopWidth=HeightCaption&Inkludera filer:FocusControlIncludeFileMasksMemo  TLabelLabel1Left� TopWidth?HeightCaption&Exkludera filer:FocusControlExcludeFileMasksMemo  TMemoIncludeFileMasksMemoLeftTop#Width� Height� AnchorsakLeftakTopakBottom Lines.StringsIncludeFileMasksMemo 
ScrollBars
ssVerticalTabOrder OnChangeControlChangeOnExitFileMasksMemoExit  TMemoExcludeFileMasksMemoLeft� Top#Width� Height� AnchorsakLeftakTopakBottom Lines.StringsExcludeFileMasksMemo 
ScrollBars
ssVerticalTabOrderOnChangeControlChangeOnExitFileMasksMemoExit   TButtonOKBtnLeft� Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeftTop�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftVTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeftYTop�WidthKHeightAnchorsakRightakBottom Caption&RensaTabOrderOnClickClearButtonClick  	TGroupBoxDirectoriesGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight CaptionKatalogmaskerTabOrder
DesignSize��   TLabelLabel2LeftTopWidth\HeightCaptionI&nkludera kataloger:FocusControlIncludeDirectoryMasksMemo  TLabelLabel4Left� TopWidth^HeightCaptionE&xkludera kataloger:FocusControlExcludeDirectoryMasksMemo  TMemoIncludeDirectoryMasksMemoLeftTop#Width� HeighthAnchorsakLeftakTopakBottom Lines.StringsIncludeDirectoryMasksMemo 
ScrollBars
ssVerticalTabOrder OnChangeControlChangeOnExitDirectoryMasksMemoExit  TMemoExcludeDirectoryMasksMemoLeft� Top#Width� HeighthAnchorsakLeftakTopakBottom Lines.StringsExcludeDirectoryMasksMemo 
ScrollBars
ssVerticalTabOrderOnChangeExcludeDirectoryMasksMemoChangeOnExitDirectoryMasksMemoExit  	TCheckBoxExcludeDirectoryAllCheckLeft� Top� Width� HeightCaption&Alla (rekursera inte)TabOrderOnClickExcludeDirectoryAllCheckClick   	TGroupBox	MaskGroupLeftTop�Width�HeightLAnchorsakLeftakTopakRightakBottom CaptionMaskTabOrder
DesignSize�L  TMemoMaskMemoLeftTopWidth�Height4TabStopAnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneLines.StringsMaskMemo 
ScrollBars
ssVerticalTabOrder    TStaticTextMaskHintTextLeft TopqWidth� Height	AlignmenttaRightJustifyAutoSizeCaptionmasktipsTabOrderTabStop	    TPF0TEditorForm
EditorFormLeft;Top� HelpType	htKeywordHelpKeyword	ui_editorBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp Caption
EditorFormClientHeight}ClientWidthaColor	clBtnFace
ParentFont		Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�                                                                        �vW����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������vW�                                                                        �vW����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������vW�                                                                        �vW����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������vW�                                                                        �vW����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������vW�                                                                        �wX����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������wX�                                                                        �xY����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xY�                                                                        �yY�������������������������������������RW^������������������������������������������������������������������������������������������������������������������������������������������yY�                                                                        �zZ�����������������������������������������*''�DHN����������������������������������������������������������������������������������������������������������������������������������zZ�                                                                        �{Z�������������������������������������}�������*''�)&&�ev���������������������������������������������������������������������������������������������������������������������������{Z�                                                                        �{[�������������������������������������ſ����������`o}������������������������������������������������������������������������������������������������������������������������������{[�                                                                        �|\�����������������������������������������Y]c��������������������������������������������������������������������������������������������������������������������������������������|\�                                                                        �}\�����������������������������������������������������������������������������V����������������������������������������������������������������������������������������������������}\�                                                                        �~]�����������������������������������������������������������������������������?���,������������������������������������������������������������������������������������������������~]�                                                                        �^�������������������������������������������������~������������������������������G���-��������������������������������������������������������������������������������������������^�                                                                        ��^��������������������������������������������������������������������n���3���F���#���L���-�����������������������������������������������������������������������������������������^�                                                                        ��_�����������������������������������������������������y�����������N���������������k���"���J���-�������������������������������������������������������������������������������������_�                                                                        ��`�����������������������������������������������������r�������k���P�������������������f���"���H���-���������������������������������������������������������������������������������`�                                                                        ��`���������������������������������������������������������<���,���)�����������������������c���"���E���,�����������������������������������������������������������������������������`�                                                                        ��a�������������������������������������������������������������0���I���1�����������������������_���!���C���,�������������������������������������������������������������������������a�                                                                        ��b�����������������������������������������������������������������2���M���5�����������������������\���!���A���,���������������������������������������������������������������������b�                                                                        ��b���������������������������������������������������������������������2���O���:�����������������������X��� ���>���,�����������������������������������������������������������������b�                                                                        ��c�������������������������������������������������������������������������1���Q���>����������������������U��� ���<���+�������������������������������������������������������������c�                                                                        ��c�����������������������������������������������������������������������������1���S���B���}�������������������Q������:���+���������������������������������������������������������c�                                                                        ��d���������������������������������������������������������������������������������0���U���F���{�������������������M������8���+�����������������������������������������������������d�                                                                        ��e�������������������������������������������������������������������������������������1���W���I���y�������������������J������5���+�������������������������������������������������e�                                                                        ��f�����������������������������������������������������������������������������������������0���Y���M���w�������������������F������3���+���������������������������������������������f�                                                                        ��f���������������������������������������������������������������������������������������������/���[���Q���u�������������������C������1���*�����������������������������������������f�                                                                        ��g�������������������������������������������������������������������������������������������������0���]���U���s���������������~���?������.���*�������������������������������������g�                                                                        ��g�����������������������������������������������������������������������������������������������������/���_���Y���q�����������{���u���;������,���*���������������������������������g�                                                                        ��h���������������������������������������������������������������������������������������������������������.���a���]���n���|���w���r���l���8������*���/�����������������������������h�                                                                        ��i�������������������������������������������������������������������������������������������������������������.���c���b���l���s���n���i���c���4������(���.�������������������������i�                                                                        ��i�����������������������������������������������������������������������������������������������������������������.���e���e���j���i���e���`���Z���1������%���.���������������������i�                                                                        ��j���������������������������������������������������������������������������������������������������������������������-���g���i���h���`���\���W���Q���-������#���.�����������������j�                                                                        ��k�������������������������������������������������������������������������������������������������������������������������-���i���m���f���W���R���N���H���*������!���.�������������k�                                                                        ��k�����������������������������������������������������������������������������������������������������������������������������-���k���q���d���N���I���E���?���&���������-���������k�                                                                        ��l���������������������������������������������������������������������������������������������������������������������������������-���l���u���b���E���@���;���5���"������6���mdZ���o�                                                                        ��m�������������������������������������������������������������������������������������������������������������������������������������,���n���y���`���;���6���1���*���7���ufY�����tdW�r\O:                                                                    ��m�����������������������������������������������������������������������������������������������������������������������������������������+���p���}���]���2���*���:���ufY�����ŷ������ubS�r\O:                                                                ��n���������������������������������������������������������������������������������������������������������������������������������������������+���r�������P���:���{m`�����ʾ��Ǻ��ŷ������ubS�r\O:                                                            ��o��������������������������������������������������������������������������������������������������������������������������������������ϼ�̬������*���f���S���wh[����������ļ�ʾ��Ǻ��ŷ������o]U�G=nO                                                        ��o���������������������������������������������������������������������������������������������������������������������������������ʪ��ßz�ßz�ßz�����?���vfY������������������ļ�ʾ��Ǻ����t�\Nl���	�:                                                    ��p���������������������������������������������������������������������������������������������������������������������������������������������������������wgZ�����ƹ���������������û���v�bTt�$%������	�:                                                ��p�������������������������������������������������������������������������������������������������������������������������������������������������������������{hZ�����ƹ��������������fYu�7<��*.�� "������	�:                                            ��q����������������������������������������������������������������������������������������������������������������������������������������������������������̹�����{hZ�����ƹ������k_u�JR��>E��4:��*.�� "�������                                        ��r������������������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿������yfX��{n�h\u�U^��S]��HQ��>E��4:��*.�� "�����P                                        ��r��������������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿���ì���r�kZ\iYLd�48��FN��T^��S\��HQ��>E��4:��&*�����$                                        ��r����������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿���ì���rԿ�f    
�M��16��FN��T^��S\��HQ��8>�����_                                            ��r������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f            
�M��16��FN��T^��JR�����_                                                ��r��������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f                    
�M��.3��;A�����_                                                    ��r����������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f                            �G�����U                                                        ��r������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f                                                                                                        ��r������������������������������������������������������������������������������������������������������������������������������ư�׿��������rԿ�f                                                                                                            ��r�����������������������������������������������������������������������������������������������������������������������������׿��������rԿ�f                                                                                                                ��r�����������������������������������������������������������������������������������������������������������������������������������rҿ�f                                                                                                                    ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���rҿ�f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���������������������������������     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��      ��      �      ?�      �      �      �      �      �      �      �     p�     ��    �?�    ���    ���    ���    ���    ?����������������������������������(   0   `          �%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�vW�                                                        �vW����������������������������������������������������������������������������������������������������������������������������������vW�                                                        �vW����������������������������������������������������������������������������������������������������������������������������������vW�                                                        �vW����������������������������������������������������������������������������������������������������������������������������������vW�                                                        �wX����������������������������������������������������������������������������������������������������������������������������������wX�                                                        �xY�����������������������������w{��������������������������������������������������������������������������������������������������xY�                                                        �yY���������������������������������)&&�:<@������������������������������������������������������������������������������������������yY�                                                        �zZ���������������������������������79=�)&&�)&&�Yfu����������������������������������������������������������������������������������zZ�                                                        �{[���������������������������������|��)&&�^hs��������������������������������������������������������������������������������������{[�                                                        �}\�������������������������������������O]j������������������������������������������������������������������������������������������}\�                                                        �~]�����������������������������������������������������������������J���K������������������������������������������������������������~]�                                                        �^�����������������������������������������u�����������������������,���;���O��������������������������������������������������������^�                                                        ��_���������������������������������������������~�����������x���K���K���2���9���O�����������������������������������������������������_�                                                        ��`���������������������������������������������o�������Y���������������Y���0���7���O�������������������������������������������������`�                                                        ��`���������������������������������������������{���a���9���g���������������V���.���6���P���������������������������������������������`�                                                        ��a�������������������������������������������������>���6���A���i���������������Q���2���5���P�����������������������������������������a�                                                        ��b�����������������������������������������������������P���=���E���i���������������M���/���3���P�������������������������������������b�                                                        ��c���������������������������������������������������������P���<���I���i���������������I���.���1���P���������������������������������c�                                                        ��d�������������������������������������������������������������P���;���M���i���������������E���,���.���P�����������������������������d�                                                        ��e�����������������������������������������������������������������P���:���Q���i���������������A���*���-���P�������������������������e�                                                        ��f���������������������������������������������������������������������P���9���U���i���������������=���(���+���P���������������������f�                                                        ��g�������������������������������������������������������������������������P���9���Y���i���������������9���&���)���P�����������������g�                                                        ��g�����������������������������������������������������������������������������P���8���]���i�������|���s���5���%���'���P�������������g�                                                        ��h���������������������������������������������������������������������������������P���7���a���i���u���p���g���0���"���$���P���������h�                                                        ��i�������������������������������������������������������������������������������������P���6���e���i���j���c���[���-���!���"���P�����l�                                                        ��j�����������������������������������������������������������������������������������������P���6���h���i���]���W���O���(������ ���@�����                                                    ��k���������������������������������������������������������������������������������������������P���5���m���i���R���J���C���%��������������                                                ��l�������������������������������������������������������������������������������������������������P���4���q���i���F���?���7��� ������ ���hd\�jU@                                            ��m�����������������������������������������������������������������������������������������������������P���4���u���i���:���2���&���"��������n`�s`R�jU@                                        ��n���������������������������������������������������������������������������������������������������������P���2���y���i���)���'�������Ǻ�������n`�iWX�33f                                    ��n�������������������������������������������������������������������������������������������������������������G���1���_���=�����������˾��Ǻ������OEx���  �                                ��o�������������������������������������������������������������������������������������������������ؿ��Ǥ��Ǥ������D���6�������������������˾������������  �                            ��p�����������������������������������������������������������������������������������������������������������������������~�m_�����������������6<��(,��������  �                        ��q������������������������������������������������������������������������������������������������������������������о��®��vf�m_���������R\��DL��6<��(,��������                        ��r��������������������������������������������������������������������������������������������������������������о��ǲ��«���p�iXX�PEx�6=��PY��R\��DL��6<��(,������                        ��r����������������������������������������������������������������������������������������������������������о��ǲ��«���rſ�j33f����:@��PY��R\��DL��&+�����]                        ��r������������������������������������������������������������������������������������������������������о��ǲ��«���rſ�j          �����9@��PZ��8?�����_                            ��r��������������������������������������������������������������������������������������������������о��ǲ��«���rſ�j                  ����� #�����_                                ��r����������������������������������������������������������������������������������������������о��ǲ��«���rſ�j                          ������]                                    ��r����������������������������������������������������������������������������������������������ǲ��¬���rſ�j                                                                                ��r����������������������������������������������������������������������������������������������ì���rſ�j                                                                                    ��r�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ�Ţ~���rſ�j                                                                                        ��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��U                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������  ������  ������  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �    �  �      �    ?  �      �      �      �      �      �      �      �      �     �     �   ?  �   �  �   ��  �  ��  �  ��  ������  ������  (   (   P          @                                                                                                                                                                                                                                                                                                                                                              �wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX�                                        �xY������������������������������������������������������������������������������������������������������������������xY�                                        �yZ������������������������������������������������������������������������������������������������������������������yZ�                                        �zZ���������������������������������w{�������������������������������������������������������������������������������zZ�                                        �{[�������������������������������������)&&�9:>����������������������������������������������������������������������{[�                                        �}\�������������������������������������8:>�*''�q��������������������������������������������������������������������}\�                                        �~]����������������������������������������n������������������������������������������������������������������������~]�                                        �^������������������������������������������������������������y���9������������������������������������������������^�                                        ��_�������������������������������������������������������������Q���Q���D���������������������������������������������_�                                        ��`���������������������������������������������u�����������^�������8���N���D�����������������������������������������`�                                        ��a�������������������������������������������������~���@���������������7���J���D�������������������������������������a�                                        ��a�������������������������������������������������/���H���I���������������4���F���D���������������������������������a�                                        ��b�����������������������������������������������������D���Y���L���������������1���B���D�����������������������������b�                                        ��c���������������������������������������������������������D���X���Q���������������0���>���D�������������������������c�                                        ��d�������������������������������������������������������������E���W���T���������������-���:���E���������������������d�                                        ��e�����������������������������������������������������������������E���V���Y���������������*���6���E�����������������e�                                        ��f���������������������������������������������������������������������E���V���\�����������u���'���2���E�������������f�                                        ��g�������������������������������������������������������������������������E���U���a���~���{���h���&���-���E���������g�                                        ��h�����������������������������������������������������������������������������E���T���e���r���k���[���#���)���E�����n�                                        ��h���������������������������������������������������������������������������������E���S���h���f���]���N���!���&���8�����                                    ��i�������������������������������������������������������������������������������������E���R���l���Y���N���?������!��������                                ��j�����������������������������������������������������������������������������������������E���R���p���M���?���2���������Yko�sYM                            ��k���������������������������������������������������������������������������������������������E���P���t���A���.���!���q�����x�s`Q�sYM                        ��l�������������������������������������������������������������������������������������������������E���P���q���(�������ʽ��Ƹ����x�THf��                    ��m�����������������������������������������������������������������������������������������������������B���C���������������ʽ�����������                ��n����������������������������������������������������������������������������������������������ʴ��ɲ��Ĳ�������w�������������;?��#&�������            ��o�����������������������������������������������������������������������������������������Ҷ��Ҷ��Ҷ��Ҷ��˯���o^���w�����_f��DL��39��"&������            ��o����������������������������������������������������������������������������������������������������������ɴ�͵��_Oh���HP��U_��DL��39������            ��p������������������������������������������������������������������������������������������������������ɴ�ּ����p�)��� ��HP��U_��05�����-            ��q��������������������������������������������������������������������������������������������������ȳ�ֽ����q���U    �����-1�����-                ��r����������������������������������������������������������������������������������������������ȳ�־����q���U            ������+                    ��r������������������������������������������������������������������������������������������ȳ�־����q���U                                                    ��r��������������������������������������������������������������������������������������ȳ�־����q���U                                                        ��r����������������������������������������������������������������������������������ȳ�־����q���U                                                            ��r���������������������������������������������������������������������������������׾����q���U                                                                ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���q���U                                                                                                                                                                                                                                                                                                                                                                                        �����   �����   �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �   ?   �      �      �      �      �      �       �       �       �       �   �   �  �   �  �   �  �   �  �   �  �   �  ?�   �����   �����   (       @          �                                                                                                                                                                                                                                                                                          �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�                                    �vW��������������������������������������������������������������������������������������vW�                                    �wX���������������������tw|��������������������������������������������������������������wX�                                    �xY�������������������������)&&�:<A������������������������������������������������������xY�                                    �zZ�������������������������;=B����������������������������������������������������������zZ�                                    �|[���������������������������������������������W����������������������������������������|[�                                    �}]��������������������������������������������;���;������������������������������������}]�                                    �^�������������������������������������w�����������H���;��������������������������������^�                                    ��_���������������������������������Z���I���������������H���:�����������������������������_�                                    ��a�������������������������������������?���u���������������H���9�������������������������a�                                    ��b�����������������������������������������?���x���������������G���8���������������������b�                                    ��c���������������������������������������������?���z���������������G���8�����������������c�                                    ��e�������������������������������������������������>���|���������������G���7�������������e�                                    ��f�����������������������������������������������������>��������������x���F���5���������f�                                    ��g���������������������������������������������������������=���������������o���F���4�����t�                                    ��h�������������������������������������������������������������=��������������f���F���/�����-                                ��j�����������������������������������������������������������������<�����������r���^���E���$�����-                            ��k���������������������������������������������������������������������<�������x���d���N���;���vj^�q`O-                        ��l�������������������������������������������������������������������������;�������g���?�����������weY�B6pB                    ��n����������������������������������������������������������������������н�����8���^�����������ɼ���������-                ��o�����������������������������������������������������������������˫��ǥ��ǥ�������te���������Ļ��38�������-            ��p������������������������������������������������������������������������������̹�Ȳ��yfZ�����]g��DL��05������            ��q��������������������������������������������������������������������������̹��«���q�YImM��5;��Yd��DL��"����            ��r����������������������������������������������������������������������̹��«���r˿�f    �+��39��4:����  �            ��r������������������������������������������������������������������̹��«���rſ�j            �+����  �                ��r��������������������������������������������������������������̹��ª���rſ�j                                                ��r�������������������������������������������������������������������rſ�j                                                    ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���rÿ�j                                                                                                                                                                                                                                                                                                                ���������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?�  �  �  �  �  �  �  �  �� �� �� �� ���������(      0          `	                                                                                                                      �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�                        �vW������������������������������������������������������������������vW�                        �wX�������������imr�~������������������������������������������������wX�                        �yZ�������������|��)&&�ew�������������������������������������������yZ�                        �{[�����������������[n��������������g��������������������������������{[�                        �~]���������������������������������>���=����������������������������~]�                        ��_���������������������t���������������C���<�������������������������_�                        ��`���������������������W���A���������������>���;���������������������`�                        ��b�������������������������>���U���������������9���:�����������������b�                        ��d�����������������������������?���X�����������q���4���9�������������d�                        ��e���������������������������������>���[�����������b���/���8���������e�                        ��g�������������������������������������>���_���z������T���*���7�����p�                        ��i�����������������������������������������=���b���n���i���E���&���/�����                    ��j���������������������������������������������=���e���d���S���7���!��������                ��l�������������������������������������������������<���i���Y���<���'���4���udW�o^M            ��n�����������������������������������������������������6���l���I���@�����������^Pe�		�        ��p���������������������������������������������������������8���W���������������!!����		�    ��q������������������������������������������������������ϼ�û���lZ���������NU��/4������    ��r��������������������������������������������������ϼ��ë���rŋoY.^Of�58��Xc��DL��%(����    ��r����������������������������������������������ϼ��«���rſ�j    		���17��BJ����  �    ��r���������������������������������������������������rſ�j            		�����  �        ��r���r���r���r���r���r���r���r���r���r���r���r���rÿ�j                                                                                                                                    ��� �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �   �   �   � @ � � �� ��� (      (          �                  �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�                �vW����������������������������������������������������������vW�                �wX�����������������hlr��������������������������������������wX�                �yZ�����������������{��gt�����������������������������������yZ�                �{[���������������������������������E������������������������{[�                �~]���������������������������������u���I��������������������~]�                ��_�������������������������E�����������l���A�����������������_�                ��`�����������������������������R���}�������^���;�������������`�                ��b���������������������������������Q���w�������O���3���������b�                ��d�������������������������������������O���q������B���,�����{�                ��e�����������������������������������������L���j���c���5���%�����K            ��g���������������������������������������������J���e���G���'���%���ibWI        ��i�������������������������������������������������I���_���5��������~q�1+~S    ��j���������������������������������������������˫������H�����������~u�����K��l����������������������������������������������������������}p�����DL��(-���鹔n�������������������������������������������������������m�E:u`��PZ��).���O��p���������������������������������������������������oŶ�m    �K���O    ��q�����������������������������������������׿����qŪ�j                        ��r���r���r���r���r���r���r���r���r���r���r���rÿ�j                                                                                                              �   �   �   �   �   �   �   �   �   �   p   0                   �  � ��� (                 @                  �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�                �wX������������������������������������������wX�                �xY���������Ľ��cgl��������������������������xY�                �zZ�������������HXi��������������������������zZ�                �|[�������������������������O����������������|[�                �}]�����������������J�����������J������������}]�                �^���������������������_�����������@��������^�                ��_�������������������������^�������o���7���t�}�                ��a�����������������������������_���z���W���.�����O            ��b���������������������������������^���a���=���#�����L        ��c���������������������������������y���a���F���/�����~�\N_[    ��e����������������������������������������W�������¶��!��
�K��f����������������������������������ν���f�te\�����mp��16����g������������������������������̻���fŪ�U    ��/4��17���<��h���h���h���h���h���h���h���h���hŪ�U            �q	�8                                                                                                                 9  ��  
KeyPreview	OldCreateOrderOnClose	FormCloseOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShowPixelsPerInch`
TextHeight TTBXDockTopDockLeft Top WidthaHeight	AllowDrag TTBXToolbarToolBarLeft Top CaptionToolBarImagesEditorImagesOptionstboShowHint ParentShowHintShowHint	TabOrder  TTBXItemTBXItem2Action
SaveAction  TTBXItemTBXItem1ActionSaveAllAction2  TTBXItem	TBXItem16ActionReloadAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem3ActionEditCopy  TTBXItemTBXItem4ActionEditCut  TTBXItemTBXItem5Action	EditPaste  TTBXItemTBXItem6Action
EditDelete  TTBXItemTBXItem7ActionEditSelectAll  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem8ActionEditUndo  TTBXItem	TBXItem17ActionEditRedo  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem9Action
FindAction  TTBXItem	TBXItem10ActionReplaceAction  TTBXItem	TBXItem11ActionFindNextAction  TTBXItem	TBXItem12ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemEncodingCaptionKodningHint   Ändra filkodningOptionstboDropdownArrow  TTBXItemDefaultEncodingActionDefaultEncodingAction	RadioItem	  TTBXItemUTF8EncodingActionUTF8EncodingAction	RadioItem	   TTBXColorItem	ColorItemActionColorActionOptionstboDropdownArrow   TTBXItem	TBXItem13ActionPreferencesAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem14Action
HelpAction    TTBXStatusBar	StatusBarLeft TopgWidthaPanelsCaptionLine: 2000/20000Size� Tag  Caption
Column: 20ViewPriorityPSize� Tag  CaptionCharacter: 132 (0x56)ViewPriorityZSize� Tag  CaptionEncoding: UTF-8 XViewPriorityZSize� Tag  ViewPriorityFStretchPrioritydTag   UseSystemFont  TActionListEditorActionsImagesEditorImages	OnExecuteEditorActionsExecuteOnUpdateEditorActionsUpdateLeft�Top8 TAction
SaveActionCaption&SparaHintSpara|Spara fil
ImageIndex SecondaryShortCuts.StringsF2 ShortCutS@  TActionSaveAllAction2CaptionSpara &allaHintSpara filer i alla editorer
ImageIndexShortCutS`  TEditCutEditCutCaption	K&lipp utHint?Klipp ut|Klipper ut vald markering och flyttar det till urklipp
ImageIndexShortCutX@  	TEditCopyEditCopyCaption&KopieraHint,Kopiera|Kopierar vald markering till urklipp
ImageIndexShortCutC@  
TEditPaste	EditPasteCaptionKl&istra inHint0   Klistra in|Klistrar in innehållet från urklipp
ImageIndexSecondaryShortCuts.Strings	Shift+InsCtrl+Shift+Ins ShortCutV@  TEditSelectAllEditSelectAllCaptionM&arkera alltHint%Markera allt|Markerar hela dokumentet
ImageIndexShortCutA@  	TEditUndoEditUndoCaption   &ÅngraHint%   Ångra|Ångrar den senaste ändringen
ImageIndexShortCutZ@  TActionEditRedoCaption   &Gör omHint&   Gör om|Gör om den senaste ändringen
ImageIndexShortCutY@  TEditDelete
EditDeleteCaption&RaderaHintRadera|Raderar vald markering
ImageIndex  TActionPreferencesActionCaption   &Inställningar...Hint5   Inställningar|Visa/ändra texteditors inställningar
ImageIndex  TAction
FindActionCaption   &Sök...Hint   Sök|Sök den valda texten
ImageIndexSecondaryShortCuts.StringsF7 ShortCutF@  TActionReplaceActionCaption   &Ersätt...Hint2   Ersätt|Ersätt den valda texten med en annan text
ImageIndex	SecondaryShortCuts.StringsCtrl+F7 ShortCutH@  TActionFindNextActionCaption   Sök &nästaHint:   Sök nästa|Sök efter nästa uppkomst av den valda texten
ImageIndex
SecondaryShortCuts.StringsShift+F7 ShortCutr  TActionGoToLineActionCaption   &Gå till radnummer...Hint/   Gå till radnummer|Gå till det valda radnumret
ImageIndexSecondaryShortCuts.StringsAlt+F8 ShortCutG@  TAction
HelpActionCaption   &HjälpHint   Hjälp editor
ImageIndex  TActionReloadActionCaption	La&dda omHintLadda om|Laddar om fil
ImageIndexSecondaryShortCuts.StringsF5 ShortCutR@  TActionDefaultEncodingActionCaptionAnsiXHint$Standard|Standard systemkodning (%s)  TActionUTF8EncodingActionCaptionUTF-8HintUTF-8|UTF-8 kodning  TActionColorActionCaption   &FärgHint   Ändra färg på editor   TPngImageListEditorImages	PngImages
BackgroundclWindowName	Save filePngImage.Data
k  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�d�B܆Ì6�hZ{��� [��q����2�����ܕ����a���/����/
���l�֭[�/
`����T��aB3^�V��;vlE5��Ӈ����!�(^1`��m��yx1���'��%k����{v��������_�� ����ph�NT�\<~(sgf�bĪ����];!^8zp���?~�%:Oރj���;��_�6��ѽ�Xۻ1|�	1`v<�7�/����~g���_~e���AD\��܉}�Xڹ2|��,�!G������<Kl Ƞ�5��$���O@5��ڙ������2�H�2tz~k���C��`1�r� � ��s�E�%�5�%�3���a�ehpz����nN����b p��!����L�w�g3H2H�_�ր�xG�F�L�  K��6B�    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data

  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  aIDATxڝ�_HSQ����6�1_�BHP �T`0g0C�Az��-,�=&����X�z0T���H/i�� ��jnˠ@!	�nbX\��d�=�3MHY��p8�?����!8�l6G��F"���B �_|����yZ�R�J�p�(~�W�������/��&,������a|���(�{�A*
����N�r�"[Ų�����*��LLLΉ�i_���ȏ��5^����CZm�u�ǥ�8�~��,o��g�z��
 �E1@`�aѽ���7���ƞBWW'X,��b0<<�]Q��~��vtfw'"0���$��U�Os������,C(���3�����&������P��4�<Ǫ��j����_����c�mj:�y���4���Sgv��;r⓺�*�5�� mjһ��n�.��~6�
#��)��Z��5�/���SP*�K4}�-���GA�8�֭����\��-zD���V�k�J������Ul�P �)Kg�BGE�D��#B&!�mK3���w(�h+�fip6�����A�{rI�hE ���	���v��&�KDP(�~�~E�_q��x钱4�QVk�3|�O�O-���    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?Cf���X�1&���Ӳþ`��e=��(�g���?���K��t���VC��w��?�,����(
>}��p��+���/�a`f�U����k�Ϫf(�u .�o��������W�+�_1��u�����������_�D��m؃-L�$���?�*��t�A����>2`�#�2�ه�I�+�Ϫg��₪i���Ʌs̬�3�}ހHhZ�vu$C�\�>��0�<g�\����Wg���oX�vMû���k�md@8���kO��;�1 �l@\����j���K~x��9LЁ��æ�g�V�A��]4 ������c@t�����i��F@������Y�����GZ3���fXP1���EA\��0�jH�*������]�&�(̊��o%â�X�D�,@	l��9Ò�x�DU���@Xښ� Ld8��h��    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd@���]�����3L߸qm���	����?�#��]@Cmذ6�3��iǪ|��c�~0扌��-���79��Ǘ���cЛ��p���Ƿ�2 `�j�kx0�ۧ�Q$�}K���cL�ݧe�}��2�	�_f��3���.�(G.?dX���1&�_`C�8�1�ytŀ�ߓf�2|��E�ӗ�W�fX���9fVw�N!���_GQ��g2ì�`��Y�b��<��/�e�r�Ê]箂p�gxq�����a���/���;/�_{
f߹���n_AQ��_*��P�������æ�g ���2<�qE�2�4�Y�����j����m�`������E�Y�fWG2T����Hk����l��]>��`[&��(�w_�0���� H��3|z�Er�x9ì�h�����j.
�b��[����a�z��o��vAU�rF\�QU��3 
+�Ed��    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  cIDATxڝ��kRQǟs�L��9u��n�~̱�ʨ�6Al1�0X��z���{�Qob� �^hED4�
!iL�9�jfM�n���{o�J��.}�p~<���s��<��8���L+߇��ӰMoD���e�A�^T�������,J0T�ǡ	b2��pݡ;��`j� �/w����O_ �H�m��t��dǵ|b�eȭf�JK��ř� ��R�84�%�T�a�T���w�C�P����/�C�'�2沞 ,��j�ˬ� �SX7?�_0�7�Zh��{�(���\�������4D��0`K�y.��|�-B��}�")�� ��:��u����uQΦS���B�+��{h��I�RA�|� Z��HwR�U >�5v��c�\���n�m� �	Կd�佥P�ߔ+�	��Q�h�]�T["fA���0�/XIF>�Xv0:<�Y�75+�M�*ȥ�Bq�p-�������F�PK,����29���F���#*���\ :�OL,��b��S"�H�U*n@��f�cK�m��%R���&�Wb����$��e(�wǾ�2{5�тZ���u�G�ZF�J�Xih�����C��_���8�9�I4��    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
y  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�KLQ�ϝ�N�@���R�����h1j���F�V���.\��n\��;I47�h(Y6PL�֐`+��R��t���̐"�������?�"B�O!	�gs�0�&^y����;�N�'{ �QBQ�����o�ļ���]	�t:��~�[|�k7P��ͧu:=�'���m �Y�Y�f��g>�LN8���N�zg4[��j���jdiD����ŝ��#@�l%A`���ø�dQ���Gs���d���y���SI�m�:ڛ�uuX�!խ��.�jj��hH&6 �����lY*k�R�"���0��i~ *��.�l�>R��Wmյ@3$6� CAQ	��Eaq!�9�0=>����.g��6˪�Y�A�`�^b3.���}��������H3��� �Rk�^<�"�^��� =�������a��[k(V�!���$P,��hx:�4���K�����P��Kkbd���ٟ%��ŮQkt]�	�U>մ�|}��ɹ*Y�S�h��l6#����Ѕ�#�5�*��"Ɋ�ɛ�1�yB�������JTj`������5/?�X�E>s̗-m�^������C�,N��]���c��a+�`���ݧ\��n'���2�P�Jx!.�w2�ov�ĕ��q>����g:v���0�qޞ�����Y����d���rb³)its����5    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�d@D�l�LYљ�7`ak
I�����%C���������́!�P3Հy�.�z°x�1�7�?��|<�����z�p5I�h�mJ����7Cq�
���2ؙh0�����ȹ[l�,��bX������0�b��_�n�����Ƞ�&����?���k�~���W�Nj=��������ÉKwn���%��o?��]��\`vZ�3�!|����y��o� �W�c�T�b�y���%d4�0�.,q��u�U�O0��3D�X�Ū&�b���+Cgq$܀����L��p��=��2�
�1��2\�������`���`1a>0;�̀�5	`���x��b7��  +!� "��p���hkU�xn�T&A �(��������e���8*��X�j���X�0��ߊf E��  O	��NV    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  JIDATx�u�{hYƿ;���S��M�*q׵�U�ڭ������u]�ڦ��c�e��������U�����J���
Q�'��R|���C-kk���mb��13��f�J������9����DY�s�
R��黦�[wp�:�1)�T+�R�C��5_���QQ�q½;gxXB����Wa��-Y�,9S���v`D y��7��~���-I��~W��Mu�j����}����X��h�d�B��{&b,�xj�4��r�/?̝�Z[�z�
��X:^cHa6����������q�D��O��A��&|����fQJ��ߎ�23L�䄖�TP�0x���A�0��&Ga�(�i?�o����i�T���D��E��TU���n4?~���q�k�*�Nd÷���_+W���̜�5���w��SX�/�l6��)�Aܼ�7����r��?K�ݻ(��.���s8T6&r�d�H���ǅ�	��<�d��$p��yQ8Z���|��EDQ��+8u�B$�ʓ���%ҹlI�`�	.�B�P�T��y�@��P�*{Η���%��U�=����<�c�r�M1Mϛ��)����Ez�o��S� �r,�s��� �,�s�F��Ȳ���݃z��O?ڨ�H`�ϋ̼� ��ǲ�e))zز-Z�o�}H1�p��dE�z��he��u�֬����F0��f�W'�^:M,�H7�CFz������@�%��򨫜�i����#����I%�?A�]����W=�T�:�`�p���$�Ƣ�>�0X�y�8%���Q���9i=�����ks����#����`E��VE�ț΍Z���Q��M?����䷆�u{ƪ{�/m�m$yL    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  FIDATx�cd�55��@��=r��u[Br���g`DR���#�AQI�aѴN�"9~I%=}C��;���P�o��B]Ë��:��f�X��!M��r`���y~��w�W�i��.`@ۗN@�>�����Ν����s��m���l��p��M����1��Z�U��2��-f��� �0l�w����o�=�ze���f���f���'܀3���V��|j?Ã��'ܺu����Fv>*�&(.�cPW�f�dcax�����/���ܻq��ک��n޼fͨ����R��B�	����*l�̷�u�4Tn�}�p��i����޽{�H���嶒�)���4ý���\9�����;w����F�R��S=U���/3�;���ë��@����q�������Dy�1�H�0\�z����S��Y4 �<ЀhP<Tҳ�s��F'X��g.���������oܸ&Ϩ�o�����<�!�������3���/]8���P�_VQ��To�{����/}-%����uz�������݃˯���Rph��h:4��<� KFP��  ,/�A�x    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd�l���Y7����M`f"#�<0����#��'� l6�h� �P�\ 0`.����R��?w�ea�|� ������+�=��Ee�J�8���$cק=:��߻���z�����a��a9k��_���_�t�w66�{K.3������������}�b�˖���R���_��+��c@???;;ûw�ﱲ�JHH�s=��0����9P�[o���yRLT����������������s;�?�X���f��&222̃1$�CU>f�bi�aaav �`�|�گ��?	>���9f���O����3@��������"7;;;�����������Ar�B6 ���h�s]c���#�������{����uG�Nf���rQk����;��9��̰�������p�
b��^��� �%�����    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
P  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڍRyH�a�}N��Gba���v977�u�QxdA�E)�H�Z៕)�����A%�`�BA���i��y�sΉό��N�����ف?xy���=���}	,C 5�WȲ���O���H�B��!yxx��$+�u	�,MOk��U#�����)�O~E�m%J/���c��׊#�b��������+�����E��;��d��w~"��"]�=BbS,��]���?p��~s�ܟ��7*��hO�x�\�7��<:����V|�(ד�Ĭ
T�_��P~��,ХjĠ�C�N�9�t�H����XnՁ����'ض���"�z;Уz�B/3�
EE�\���a���Aؠ��:����Z ��r�<���+�_��z��j�ϙ�z}w?÷�4��i15kB�Y9>�_�RQ#U*]�|S؎Ί����#�Y���IH|ɛ����kj�e�ɉY��zH����E^�Ը�<))�=���e�WJlB:��nF{w?�rN�x�[�~b��r��ñ�7Ρ��=$�3/GL��4�;*:�~*�@YA�����`gk�-�|�>,�
��0�#�e����Y'�JZm���3.P;80_U;0�q2?��Ъ���%sCU��FF���,w�D8��O@�F�8�۝�.Q��nƇ�X'|��AaEP)��x�J��4&�����    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  5IDATx�c���?%���ѻ�d�PH���F�?ï?ę�7a�i����,`(�u���D;��~�
���30����\��g��� �o?���	��700b�y�:� �7����-ˎ��g�PԿb����/��ܾ����S��pWc)��OX�0����������G�Neؼ'�f�/J��bwAi����$A���F>��[�}�W'��,�l@̺�@�@�`��i߬�h�w_��+Q�Al���j���"��(Ԋ�݀�@b�|!�U��Q���Gz^�87Rj  ���qx    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�mSKLQ=3�ϔ��P@
���E���2��Ѱ�HPQ�G�l\�V?$�� @4ą���L�5�������Ng|�P�[����s�}��m��a��Pb�@�E���R�GA�^:^��m�S�^*��!V�H�Ȯf��Ӛt�JV�b\��+K�;5���@}4!�yx4]�U�k*��n�!��x�J�,��<5p�M"��|$"5�"�@Q��3��p�XX&e��&q�5MЪ�fx0`âXF&���A���l_���4X�@i-,�G�4�d�w\���\�_��ǣ�@P�1��A�pL|#;WA��gd�鳌RvK�m[��a�~�%d5��=]���.�M�Uz�Xq�w�ak�y�E�Tm�*i�̡t|����tϠ�V%,Ez\x���RL�E�0���(���x�����p��b��d���2����H*sLI;-��tX��#&���1�՟�������r�wY�
6E�EKX��nG
�F��0c�.Q��n��)�l��d��çb!�����T#-*��(��6�ͅA+Gs�\J�����
�H�s�]JV}Y��#��~ތ��]SIq��"��j����J�ʫ����M���d��*ebo/��ꘚ�&��Qɟ�íl��^���$L����#kA����ñ�I?��U�8����VJD�4m��D
�d��3�w��V�_l�'|=&.    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  nIDATxڍ�]H�Q��6Ge6����,���E؅Q�2�ӥ�H7eN3�ۖ���.b4}3��o�&]ɊP�>�p�+A��s�6���A��P��꜇���s8�p!(��!X58ܵ�$ma�38�e���5/�㢳�x�w�5��o�z=2���0�J�s�+>ע��9]�|�����!��I���pY�Mt�,�}+Qkx��]���m�Ö:YJ�Uv�����g�E��_V��$��~	<�1��+!�$����R�.Ut����܇��F$=&��a{��.���[�����M�,���6r=�����gڶ͎��"��L�/r�4���@���з�1��]rv�[�?���B;�՝h��Y@B].��<T��I�,�C��`�ly���[V��X�£�%]�ֶ�"�2�� q73Eg�2Qt���WzK݊f��2ʞ���, �چ��-�ݸ��y����X��d��"�ĥ��� A-���#0O�<_�ߑ�-b�����#��M��t��R��%4��rq�D!�p�f�z�N��G|�.���N��O�:����Z��i�z����>�Y�S�
 m��p�V��?�.�w�    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  [IDATx�c���?###6�ట���?�b*��D��`g����%�ψb@C��=��`6���s������L����3K�0�?����o�H�����+;�VAa;e~A���/_�<y�������hj��\�r���� Fb7l����PV�d���û�����3��3���3�}��P\RZ����]�(Į����ݢgd�����;7/�����F�(eu1q)x8�<�� ������x���^8�����&��]U��,����IEM	Aa1��N�G3 n�{M+���^3<}t{��Łq I���Kɫh�J����31��a`����]�����?X4	b���@�#~O�_�o�l�W%MS�o_0�}���ᒀ2 �)6�R�`ffex����?̺����!� ��Ŝ�<=�@�~����0����`i�	�\�����_�˼|B*\<?|c���=ÿ��n����)P��K�vc5 ���+���p���[���,����!���2�#�_�{��na5 ����gf������&ffPB˃\4��ޢ�=8���LL�@%6@y -T�Y�`,w�@	  �7�_�!W    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
E  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c��]����������Ł��b�
���{{�2��|���?���b�C����;vlex�8�� OO�NTqP��/��]۰������߀����ف� 7/�f_�xƄ��#&H�a6��œ!߉�A�����`)a6��ك��?`SO��@J���utg�5��ѽ��	� k{7��?!�;��9Lp��u��	1���n��S��x����k���w10S�A�d%MFFF�+g28 ��%| ^@w60����2�a�a���ã�a2;��A�����w�}aȜ��AD\
^X@�9V՗4h2|���#��d�����0K�Q� ���<A��K�˕>CH���ATB^X�
5L�U^a��xGL��2 �r���    IEND�B`�  Left(Top8Bitmap
      TTBXPopupMenuEditorPopupImagesEditorImagesOptionstboShowHint Left�Top�  TTBXItemUndo1ActionEditUndo  TTBXItem	TBXItem18ActionEditRedo  TTBXSeparatorItemN1  TTBXItemCut1ActionEditCut  TTBXItemCopy1ActionEditCopy  TTBXItemPaste1Action	EditPaste  TTBXItemDelete1Action
EditDelete  TTBXSeparatorItemN2  TTBXItem
SelectAll1ActionEditSelectAll  TTBXSeparatorItemN3  TTBXItemFind1Action
FindAction  TTBXItemReplace1ActionReplaceAction  TTBXItem	Findnext1ActionFindNextAction  TTBXItemGotolinenumber1ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem15ActionPreferencesAction   TPngImageListEditorImages120HeightWidth	PngImages
BackgroundclWindowName	Save filePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  OIDATxڭ�Mh�`���V�@�v2����
T�u��֮�hq-x�T�"�'A�2(;)���t�ã��V;�йYR6ċE���#I���m1s�<��<�x^�T*a#�������p�?�ė'΃l�L��>�b�K(�"�Ţ�D��"�ܓF�/�&p-U�nw���
~��4V��/!�A��!/b��&p�y��pPZ�2X��6��h�L�Ԡ�j'0��^+��H)���ݖ^���:iM��q��X4��=��ry���ޜ,��3SH���lEF/v�h��oX�FBe�]lZ��H�M�)cn6V	v�,`��޾R����n0>U��{�����=M�7QHg9d*+'g�5�}�hַV��g���n��\��w�߈c�=�;y�8������3��*�i!�� O�XI����0�J`GK��_�q�5�K����,�U"���30iN�6<=��r�t�6�6��a�&���I�KeP(��<�^��ѿ���z���l	.�Wr�sѠi��2a��7lW��J��(�u�y7��j���w �ק:���}��=Lm�/�'J}v�ƒ�    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  %IDATxڥ�HSQ�ϝ���4$F���ʢBgE�"��Y��0�
���mE��ֶ,�Y�Qն�)�i��H�,���D,K�m{�������Қu�qx�������>~Zvv�I���ժSƋc�}�ۼ9o����^�l6�HD迁�t'N�>%�h� U��dd�,�ٚ�4]~����]�ri�J�"����̼⸸�-K�N�I���t_�Z?[.W�X\�x<^`hh�y� /�Á���:����@�pח�ZE�R����bMWWTJ�����ʪ���O�z���7�����Jk���Cױc����L6��o]����'�/��hGdcc#TT����_��fX뤻,lu�Z��ܶ� >4�Z��q:�YOF��L��d�� C.FKB/Ix1}E[�9�r��1�zSs󭾟7��9�ڊ�@Kh쾏 �Hx��}L�
���@�
��nk{���1�kc�,n� F��v$C{�����\�i���ۃ�7�A���2���p���7��\nLﶛ�7F⌰���Yq�����!!�iK7��x�X����!�>loW���tYQa�T�Ya����TAS���.[)eR\���,m���Dwr�M�N�r�u�0~� q��ǽ���|�7�L	�����2��i7+r'�2/���������R���q�G��)��@�_�M�ґ�o'��f�̉����k��@��T&:�0�9�$%!�,,$)&�W�������_,aw8�5��h���������������IXCdLc��B3��|)~�rY!    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  KIDATxڍ�MOQ�߉��������X�)R���p�G���"A�i�-�i-
�P���$��Tх��IZ+�u���#6N���.n&�s�99O�p�\qO0�ͧ���ɱ�*,�r\�;E|7N����[y�je���|&_dB��Kw&ɠ�J�7�p+�`u}c��.BQZ�"�b/L����/v�G��i��|y��*YNd��IhGV�E�py-��_��k�/XOsL���q"Y5�)�'���2U����{���w�u��7Bd�������{
��٥8&���eՁ]�p��,�'���`7Y�xљ�7�R81أKU�q���zB�o�#+��
}�7�6W���D��x�j�L�������?%�d���;CDvvb#[R5��Ǡ�j̱�x2���MS�m��`ͩ
3�h��/���BС�y!H$�������;��ƘuG`�Dr�5��"�hDbS��}�,*�3�!Q_j��o��ih�sMs�{�]gk@���$��!�,Z�(�{l oRe5�j�!�<a���cu� U-w�~#X�-M-N�0Fow��gL~�+�D.p � ��4��    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  dIDATxڍ��ORq��O/\smݶ66��n���LAD#AK/2{]��(���Mq�V�"��T�tԺ�e��5'!�6L%E�`���I����|�Ϟ���0!�ZB��5-�\���[�=*�Pqk;P$*�;� �E��*v���s)����� 8�h�5����Mb���᳃�ٌ����r�Qo�P����91�	�Nj�<dG���R,x���i��v!500�θS���?���N�"�[����`�3N��Y��
,�D
,I����1��B�I^-���Û7z�}��Z���n��������u�5� �C�~�u�`�$�H��U� 	��pPC��W�Q�����M�GfF:|K!���C�(�� ��"L��)в��2��ש�и6�\���=���$��B|wب��ah����lu0��}�hWI�`^�	L�G�p���*���5V0�B��
SKy��/��6L�{�\��Y
��-+���AkA�Z���x�韧¯��`h�a1Ⱦa�v㑦"fd�v����0�+�db���$ʻ�𸭊�l�*�;CK*�O�yC�ʚL�^-�%�#�Қ�u�47(mlg�b�oU���[l�L��    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  iIDATxڭ�KLQ�ϼJ��T(�vڢ�� `�D0�F�#EA
�w.�jĽ{L�,�S1Fc�h����
ʣ-�P���ii;ӹ^[E��$��s���?��g��� �@b[ͮ.���l5߉*/��*�D���8�@���/þ�@�![N�V3$���V:��XKщ�$ES��,e�Z4EC(�i�<�O�Ũx��v��@��s��e��V���3��\��5V�k�$ɟ>�����wo�����Z�����٘�6�Rf�p�<hҵ����qO��)�C�J�
c�}�z�~��q��X�5�䗜^���?�8G�`�#w��9 a��LQ�YSκ�4M�}^��mwX��mWr�66|SI���׃�A~;nxϧ״+�ɲ��e�Ir���E����Vs	����ɺ��
�f��$�`Ň|��ځ�x^_gۑ��y_o���8p��F��|e^��т�
�b�0f�����VY�X�<C���4�[�I�g`t�u�X˾�	`vc�G��ՈBD�*"��Q!2F ��	IB��۪o��!k���J��CA�ms�T�%���#_"�t@��8ǣ#�?M���m�)�T���o�j><?)�W#f��Y����4#� ���0�v��
��0k��dF�}�ՙ6�dr��rA��R�n�k [�n�\T�i+�T1|�t=vX��.��/�5�U$m`h��H�� b7E3�J�
��%�\�����\�����[���f9E1�h�I&(�c�P4���Ql'�(�b��jUW�fK��RUK��|��uż��x��zg���?�vI ��)<5g��b	Ũ$��f��]Xl�?����D��ʋY#H{��ډ�.l��W4��,���    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  CIDATxڭ�KLQ��<:�N��R���#"!Qy)�R��ua���VM�,���Ġ�Ld�+]�0!�rS����>P�
HDD��Cg�i�3�)O�ݽ���s��/��<�O�D AҢ�t� F����=��^�U��nA<t��I�$P���r���"����@������;��,mjuVGQi4>�:T�q��H�*ӹ\#>�VT楥�A�����{��P���Ͱ���M����# ���1w���2��wNV�,uJ�j�Py%#�D�C`r|�G�$�^o��ך-O5�����Àe�`��H4�Oo)���tYN��J@QT&E���@(���� ,���9y�E��`zb��)��i���)@�/�V+���-,.'d&텂~�{fr@x��N�o���J��E<M�-����d+� �����PLf7��p\.�-%u�VZ��L����8��6�v[�hG��+�ޯ�/��r"�l��/@�������kG��L6�d�4\?��8��8l�ۍҮ�ާ���8�H9��E��������T��-3K�Ae�zf���H�����RW���k,g}�����<2Q��%��E���VB��]��X����XSo����NU�Fð��1�$��#~�~u�^)��$4���������'Xkn<���Ge�Jf�`YQ-�\�:�Q)5f�s�_[-���'��)J������ 0�H*�������N�5��G(��G��x���ŕ���K>V�X$��0*6��5����os��'��������~�d�"�����}.��a�#�B<��q�U��۵^�~ھ�u�����:�    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  CIDATx�c���?5#�����T1uEg*#����)_=��-��P3���h~���aݞ��n=ax��XL���AWU�!�̈́���E}"��������m�f�G��bu��� CSv 33\,����M����x�Q0[_]���P���.0��qmE����8\Or��s����^�c�~�óWb},XX����O]gX��8����`��דR?��YH"���1<}�����'/ޅCr�=���2\]��3P�q�9Þ�Wn ]���_���PLo@3pF=��S��2�[w�fzWCQ�A]Q����_[]�x1ؑ����hN�O�K6O� ��`�곃�x�����fX����(f6�G5pZ���� q~^.���pFF����N_�Iw@/��(��d5�8�a`��u/�|����Ud.�|�p����/+[cu$G�8���W�1,\#"�5�.�xf��0�����r��\����������DyLu���<r����_l���p��-P�X��@	�oE3pBe��H�iP 7��  J�I�^�D+    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  rIDATxڍTkPTe~�.�eY.K⅋`��4R"%ָHt���:j98��8E0:3�P���t�j�`D	���ea1�˲�.{���3f��g��|g��<��\ޗ�=�\U���h���[�QW���yf�M�꽠 ���u��\nm��s��Ωն�l**��C��p��@(,]��Q��q}zP]ׄ+|�35>bo.f�8�QW���j�֤m-�[�C�5�깆W�HN\���Å)�4Z�D��n�\,|4%	�wva�0U�����RCSm�|�j�T��;Z_���Ƹ�(�@� �b�0�P�݁�ch�ЮoVW-���*)�Y�QY������G{��| A2?8ICô	f�!� x<��|[;���o�4T�ϯ�p��@�|����ѭ��Ͽ�Dz�D���J����fǜ��׃��Z/��.s����ۀ�*�)/��rq\�245�ņ'W��p���z�T���'����Nu���V�A��l�1|ʹϐv�b�oaj�J���g��;��Q���p\s�ݹ�2�2T<��"��!<4��L����.�ON:=nO#�=vh/,<~n�F�"���4�08<�\KC�w�t~-2BQ�����@��Ho��,�%AE�Ax��
��,�5Y�q�"�v��-?��^}Ssc��V^Q("K}r%s862�At�G�5 ��o��Ҽ�+�����Џ�p:�G���q�\�Q�!����0ի�W)EF`YT8ܤ��j��_.�p6��oJ��C `�֭Iߒ�P<FF'���wwH�!=� 1�K���Y_�%'�xݗ��lk�g�����u�۱�PP-�>���y��Y��b��X��ÿX��q����ž��0�L���ڛ�r�,*٪�����;@ �:q��eQL&���j�2Nz[x����}����ʦ��RT:���P�ey��9O�3���H�k�U,�*%b1�S�H�����z4�"_���Ew������X�??	X�/D�|�n�7!�ν��Ɖ�OӀ�\��P��n�� ���>��u�aD;b�.ޒ���璋Qߠ��c�VX������}�����=�S����`ְ��7�!>�{�3����Ca�B����i���{i���X�	��E'    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
_  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڽ�mL[e��׌��m�Qfd,}�m]��� ��1'nat�St�D�/�����Kbb�e~��_�f:��8uDq2`P*}�-T�z{[��wұ��Q~p�'�y�}�/��s��RXR��Yj�l��l��%��di�;�0�l�rrs�����������u�Dp��H�LyMc�������8���p��W��(���K�ax�!\�܍�n_d^~��ޙS��'���M�7ʺ��7-

�ܼ����+ľ�c˞�>�\	�-,��HVJ���۸I�W��t�����va:�G8�@���z8]��ڋ��Lh	w��a�X_��7���t8l_Sd.m[J�W�7�g�)z|4�&y��SR��l�����jm��y��J��Ï/.�:-�X�E���A�w�J�"Ey�`�Z���k������cRk�S���$"��aR����8M^H�3�ħ��6���83cm֬�T��ZU�݅��,��z/>��8��;�t�H�z��R������17/t��^R�dǚ��ۺ�����`�H��n�󜊦�_�B���9��C�i��v�bѽv��J,�=��qӅ��GQ�Q��	,@,2z�&���9����X,o����}�S\��"��&M�\'i�z&9�s����s�Tn�0f# ���6�l���ͯI$�����}��4�;i����%2ç�������^��$%B��;�p6㞀�4t��:��/�R��=M�4.�w�>�o"�%��5M��vբ�P�Q�˒�p��Y�ׂ���xYuCi�nw7�E`��Z���\j�������_���ǌ���
���EZ��X�5򨖶�	��{kU�����nܾ`�z��菞�W��Mr�Z�.hj�F���<h��7_�;��a�|��\���Mr���� Դ<�
��X�؀5켵�"�ߏdY�91��Ҽ�    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATxڽ�mlSUǟs�ۗ�])[eLْQL@��- Q4�lq��mp[V�5?b4Eb����`$&�ގ%����n�ӌU�F@�c�4[��������∸��or�9������x����d�,CB�x.�_�-&yZf��J/�w��E��60
y �{�<��r���]N5ʓ8]��Xr�˻�g�`
�` 'v���y��>��jG�8T��8J�۝[@�bR�@K�B�׆x���������϶�4���V�2�
--���O�wE�Й;,U>"���=�h�D�
��%@s��	�3��ÄA�;N����E ��fo_�ͬO���}O��hn�� @G��/�����&���9crͶ�5�$��E���u��R�{�K�WpW�(�����_;[���z�N������ڌ�
�]ƨ ���2F� �EԞ���������T��8r�/�Ѕ�BOa�#{@�*�"I P�Zp�\bb�������)m�0�Z�x�7p��|I#���#"�_��4���4�&���D"	����hΦbSѶ[��'_:��g��Q2Z�*5D�Q`訲�R����8����#���5��� ��H���D1���B�;Y� ��i�_�(z�Je�V��p��op;��R��n=Job�Xp�7Ȼ��5��%'�=��+j�V$�k1y�
�=U݅����߅C�yp�o���t����pܸ&4����	�ݶH�h`m�tu(,�u䩖��]o�i4y�)p;��1_�ﯓ�J�sD�cĂ͡�:���OO���Q�-e��Q#Y��Fa��h����!��P(t=�N�R''����C���FcX?����Gϼa��~�5]�$(�GI=��R������S�/��W�Ɍ���6S9UϽ�ϩ��*�p�ک�ǂ��O��h:u�=X��[V?"�A��hkQ�8�at�+\:VS�-߅)�M0}ǤT��eDڛh��TPN~��(��;��I��ݿ���͸>��~�:��O���DBU�]    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڽ�kL�g��o��Q�f��Z(m�BVaDN�%�̒�u��:��nY�i�FƖ���x��/ f#�MZWj��Rz��YV�XZ���DP��>�$o��=�<����X$,��\J�f��l��"��>2Gtf���܄j�ǀ��W��`d�_��iP�������nK�J�&�������Z�����O�EZ?~�$��q��؋o>�-���~���ʈ��l�~��:t���k�O/ i4ZRJJ� A �HM�|���������p���`2ٛ��Ҕ�;�D�(7�f8vL�y09�c%��a�{q�K����I��_4��c>w�j���Z͗�.Ҵ�������ˢE���!��G�ݲ�]���P���߽\z8z����f���<g�H �*G ���>,���HGB<N�N�7�6�^��u��]��2B!�2��!��f�@*��wttB���h�#��d�R�N�'��n��R��\F옚�#0��f��V�l���+W:WQ㧃dU4������n 3�s�v��EF�ͣ�H�UQ�;�D�U��o���q4��|���Gff��g�s6��D^A!,F=$E���OB������]=2b�����ٳ*y��-�Q)*�r`�+)(pA��Q�75�?hn�j������l��|8ð�	�+_�	��)�\���ש�/ʷJހ /��fl//�g?:`p�,[�(�GA���׃!����G!2�c�C�WVl�3�z+v�l�����ء��c�?�źp8�V�˥�}����n�\��4h6�׈ ��ف.�CC���^�Rs�|��/�T)�n�e&����5D��@D,.Gu,F:{�C`��<.Z<.��5�~]�ʪ��K�BM����w���ݓ�N^��_�Y�~�ET����C�%��b����0��$�&JA�y��t.�g�����W4����^���o2i�0��>�    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
y  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?5#�@f�&�l�00�g����~���nn��͘�wm�?�ԟ�����ePk��.������u�g�2|���dL���(�~/��?��?Yr)�c��Y�A_�c�[H���!.,����Q!v�=�׮����W�������_~�%مE0]ݽ����p��E���^3lj�`��fch\|�(��cm��G���������cxx�6CM�6���I.,���@(~��	��+��O � �/�tI�ZL>|p�����e�Z�$������~3\�x��ח�[��9�:�%ʠ�HkT���]����M��_���D1�����X.�_40f�A`����7���3q���Ϯ�fx��C�J�\XqaE�J̜[�����7_~����>,��,6��1�*���������g�ő�ª��FUͣ�<�z�Mm��U�w�    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
X  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�}�]L[e��眞�~��t-��.���+�f����hbb�%BظY�3s��&�Ll�k��̌�F�9��c��RJ�~�����7��|�N������y��<��s�:�s��`���vP?ì�P���P��<nMV�C�zG�����򤹥z�:^�g�r	�\�T�l�QUQG����N��������� @�K-j�
^a����,���Q���L��j��\$ٌ;<O��t�* ]Fzs]O�`5�XI�̩px�Bo0CQ*�hY���.����ˢ�����0�Rkx�)���~t�$�S�-�܎�����#O

�,�E�T�g|sm�k��!O�Wo4�>�[��ʙc���?E�3
���f���bg�mA�����bu��i����,7�2��԰�3~�����)�k7ȸq�0����h��>\ ������h�p��k���a��.���b�l�Q*���#������+�X�˻�lzk��	0�����h�k��IbOWh�K� ���,��^��w�����r	�����{$�uy�L�(�g�dӣ��}Ȍ`����1$2�3]%c~t7O�ή��8�/w��~E:�4h4`d�^�������ya_�����N}D4Yn���e�V.Ѧ��vL�}�W��$�V�۟G����H&V��c#Jƛ�]M�������s(�� RS�f<�b~�$��YlvW� 6������=y�M�KJnX0d
�H���`�|��z������9Q�����G!����C�l���LDP��C���������$��1��� ��xK���ֺ�ᇡߨ�Y_�����3[[Q?����vfS�����_����LC�{�<�a�1t̲�NF
*��9�\\&N��}�7�iz��o���8��������I���T������)�>�?>����x    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  /IDATxڭ�}LMa��u�^�a����ͼ�4����P�y��ܼ�e)�sQI�4�����5����2��nuk�S�s����C�gQc~ggg�y������{$��ϐ�����6����/b{z�VB��.��h�S����~���giY΄������������Fiu=�:����1���w)�IJ�2���_���u�,u,������H�\�B�;�=$�w�����p5w6�^j���☽����8v(X]VS.�Q`x��ܽ�]&��#��i��֢��l �:M��k0��)`>E�˜!����!WB�aI��2�m�&��-w�`��.����C��J!`��~ ab	�8#�5�`"<ipۙ�DzA'�{#�=nc�ٶ]�1LE$�D�p��*��<3!5ʋCO�#���ha��u7cĠQԿ�ҽB̋ ����Ҽ���\lj.�[K�!'�j�:4w{w��a�0�l[����r/��\:��7�%�h�߂�E�2�1>4|$��X�ވ�7���̼Y�-�3ˑ� �L�xWc}i0H�MT7����Y"d@;�q����4�B��p�q.�/�!#ޏ�U���=�)��
�. tZ<�N��� �+�)��$�;x>�4�(���I�����:�m��J��'a��i�o���kC�8vs�����i�����n@#6i�"j:�j�k��D��^�ed�L�F�{��m+Rn ��&�}�0qA"�5|��l	m-x��C�A*��j�"97�Р��KD�?ErrN���Z�%z�o�裒�d    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  [IDATxڭ�YLQ���tf�QJ�Ph��FAE�"4&�DB1j�������>i�Q�L�OL��U��t�,RYZ,�zGmR�x����=�7�{�A�,��\(De��K��oe�=^��;����ӱ��Y_`�,�~	�Fn���֢��@�:�����C42�	��oണ���d2� �$9:w1m[�Y@��_�7�n�ϫ ���,�%I&����NGW�k��L?Dفlkݽi��Ǝ�z��e�{���(��e>F!�� �N�E60嘿�ǆ�>�z=D#,0�}Ma���i@G��c~��9f|w��/E	#Y|"�� t�js�+u�u��#1x�9�Tw2t4u�4����WA
{���aOr�_>ܾ#���s,7���F�� ��q�υ�u�3@����s֙��PFb��"��w2�p��4�UT�ZrZ^9n
�/�`.m^��vu]�5�z��`�7����� ǥ����zS�Sf4Y���iU�^?���\�2G���*w7�:���W��n����_�_k0ǆ%I�(��ӒhIFG��������o/��p��1-�~���:�n���4�0����V��;O��y�2���W���g�v
K�tL����%�M�04�8��W��쯀J�q؏gX5J^&c0�����WvF���_D�d�%ߪU�9.��ς(~��낄zeQ�JB�W�g��fg���8����`y��I �|���������ر�e��)5ʙjl*���D�=L��l�=�O�1i�6OD�;�����c�z7�����@FyXʰ�-�N�����ר���	    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c��]�����D�����$�eB�o?��
3�x�$��`T�]�����y��1ÿ�����@�/���lc3[��͛71<XȈ�@//0gB(3>P��/�޶m~�ܽ�������k�6�:�x�9]A�,[1pߞ���sts��X�b��;�he�
�T{�0p�B$�&�`���=�MJ�4�v�����=��>�@#K'���@N��7s�K.M�g�fcdP���@N��6��Kn�`0(8����krbl���-\r}�Y�i�/�0�����|FXL�XTJ,�,�����"�@l��~�f`h���>vh7�T�2V���De�Wy��xG�[������KW������@l����o��~1� ��>�d��|�ANI�������JZs��a��7�а��b p��A�b�}iM�a�.��3�)Xn^8��@\��<���u CS�&�@\��@��E� �#,	�^j�    IEND�B`�  Left(Top� Bitmap
      TPngImageListEditorImages144HeightWidth	PngImages
BackgroundclWindowName	Save filePngImage.Data
P  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڽ�KHq�︹�ERVf�C�AE�k����n+�%�A��D����R���A�T�S|���eR�(a�H�ή�3��h����C5f?X~����gf�aE�J�߀ކ7����=��Ҳ#@��A9�vC�~��v	�$���rx<;����ddef����������@^�*J���2t��p��--͘(@nnDQ��&C@�c����:�r�BI�:��P�D$����8� ���p�i��l��� �<�p�.tw����@�#A^���{p�>|z���=;.�2�1�Jc��� � 6�3*p.̈́�u>��׽�t #�	P0t��5��H�9�,|��X3`g�eC�t �h6��s@�w-㢠��8�蟠�y��g& E��IƆ����>���ӳ0��"��'�`�6mފjO�5����5����,Y���`/|"H��1��ϋ��xX�ccb2ʝ���s$آRxo���5<�?8tĎ	6�X>��9n~V/A2��&��l�&�:Rp�Y�k�K ~����I����Đ��ꯈWJS��d2E.���*�Ⱥ^�4`����bYS�%e7��1d��I���'W̝|>b�>�{�al;UW�B��9���?�[6�&,�z��2�,xe�T�8�f��c��    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڵ�}LSW��m��R�l+��b�,K�$-�cs
1c���Mp[����uqTܘn18C�:2��\��[ �_mun��aZ>$���B�ޝgé��N�r��=���9��C(�@�G����j X]];��W�8 �!)F�]{�����nUCC��$$$}���w�����H>���Uܱcy���s �C%������ʁ�$&&9
���9t@��0j��ǵZmZ� ��������e������ٟ� �S"S���嵸�XHO�������������� ���(���cZ�Y�����H={�ʲ�; �O�������ۛ�P(
�\�����'�������_� (..���R	 �e��,��g�smnjj[@���0���>����вN�����m[kk�w�vN��e�
P����
�]||��K���;R!6v#\�x��� ��bY���7;���ݯJ$�\T��5�D�җ��j^���v��l6[	���Nz��w�}P��d��v P��M�"S`1�Ii�4�i���w6B]]vP��M�Q[[Q��r����(\B��	Ы�!_<t�L�l��"7�ׅ3��� 5tuu�� ��Bm*�"��V��89�$�_Q�#~~v5tڪ��rEX���u<��G�'|%����25�����o����*�B�����j�𷹝��𾵛�v����[�1�����}5��9���e��=0��%c�H�uJ�@��k&��}>"�6}�zfe�R�������,��;�(��~���ׇdzc!�J�k�p��`ܾI� k���䄗��B��Y#B��Xy�yۜ]��#��B�)%W�;\���l����{F��-��i�\�V`�H����'2��;���ձ���M,��	 ���i���X���6�~� ���@D�8��x����Q�:1�%����f+#�-���*t��P��P��>�g����D�J9G�}:[a|�����_�?��N���    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  cIDATxڵ��KSaƯ�9����HӅ%��Vi���LԚn.�*�����.LT����DT*�����^�f{s�W��6\c휝�������s��P�ld����)
5I�J��l�����,���leR��=������'ً,|^���f?��g���'˼���'�|7"�5���hΟ~|Yb����#/��������se�w2��q��G$������7��0E�MUX�$9֘٥�*�i�"��S=�WY��9�a�/\�^*/"	��%��Wǉ����D��?�eX& Դ,@�m'Ɩ������<�8��f��zӀ�ˣ�n=�%�H��a�?zA�9\���4���0��ka����|L�fL��p���+*�4���1]��'�� �m����{�*8�q��*	�'ް6�����i����u
�����|1u�;X��?���>�i��0O��R�Ե�$tg�!��3p��q�v�o<����?@��M���˴���1���d U���T;�iZn��@c�æ�H����G�;���?�^e�4-7�vmC�a����u�8M�O�~�W�j[����G��H�	a ^�s�ld�����Qh�;    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx���[HSq��ꡐJ�"�+�4o���M���dI"�]̴����R�
��Y�l�S�)��x�{j�>�w�t����]��~{8�����}��v��EQ�
�P$���=I�][[�
�Sok �����KK�Z� g�F��J�Z�g@(z0����B�%�I�'�2�2�+���m��n�๱Q�|�t�����>hO�E4&U{�.�1���Ks��[������<�T�m�E�mk�z`I/�)� [�0m�����虁k��zh�I��G���GE`V�o�Y��TG�Fz��dߥ-�d4��8�t�:ԹH�0ч�<p����_{���5&�E�.�cf��X����֭$ڇ�1:����V2Bpi���&�'b�gg!��x���`�
�V���������:I��&�!���n@G��U��� �n��I;Mϣ�{�b�j
��M�'\�Ɂn+�*�0%K��ͧl$���:r�/�]2ނ0L�wq�ҫP�d@v����-��!'!.���&��c���:�?ũ̭��ؐ�ԡ$M`��y�����{�/�i�״�m聬'*�eD�/�n�oa=�{S!O��v���Yr%���,��P�vY�p���h��~��\����<ˊ1�!!���Y`�P�Ef,4��M�-����83p��Q,h4��F��e@.�C��6����'�ST�����x3��:k���1�K�Ypl���J���@Q��UXFtz#�^ƌ�oQnA�\��Pg�`�����E�    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  +IDATxڵ�_L[U��so�_ZZi{�AG�2�F���dӂ�,��e/Ɨ=�`4���f�Ąl�Z#F�BF�f؀1���Z��@{��?�[G�B��NrsϹߟ��}�;�"Q�i$B�����[�	�x/wXǻ�����D�(
S��h[x�\rW��r7��\ BV��w
D�� D`�1�X �tXYY��4_]Yc����΂@��J�i3[h0�@�����f3���`��d25�"�'2�=�ri��\�V�a~�6��bc�@-5�Z�d��e,�ϻ~��Y���S��(�����k�?2>k��0?��t:}�Y"�D|C��D�8#�8��bн�-a���%gb���\{��D���|_��T�����%�~�KMФTiް�ց��� ���@4�����X�'�j�jM����ܭ)�x�fp��WؕY�=�2��s�T��8���&x.����g�{3�i|�YC����w!]��	μ����n�i5U2Z�«9?����|�|�/�t��)(�����ޥ9Hl�������r��)[m�k��r�o���47�t���\�T��cu/xp������'�\zX��?_^Qu��z��4,����8y���9Mi��F�Q��i�2���z��kɈ�s�K �g������u�U�/�Fۏ�]�� @y��s�V(忊Rw�b aA���(dX�Hg�Xv�n��Z��wsu}n�4;Y8�=�JTZf�x�Қ+%�x��D�8=�FsM���B*���r�&@;��S����z��lom~�8�:4@rN�o�T�H&���p��)��Wڣ����
�B~
_��e
�)�����9Q|-,����_�wU��~�h2� �"@Xӎ[�Q�PPJu	(TصLn�q�����̛�i"�t���V)B� �5B��}�;�l:}#�'τ��b��	�9<zС�D_.�q\2,�g�(��o�c�a��3h�Y�/FJ�� �"��x���U������?�����h�}�D���|k�`�;B�,��#:�9�
 Os��B�۫�    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  :IDATxڵ�]L[eǟ�ٞ��Z��n|�-s�4���3���`+K������1~$��hTvc��E���b���
�B"-H�P��:aA���ў��sN��}�v���]�ܽ�����9���C��iD@Da������w-�����?ݡ�f�
_��q�-�V_��2}����I�3I?J�V���i���Q\c2<Կ��s抾#O������gqXL,������o�F�ç��I����(e�S�P� �������w�[�f��ݜ����o'¡�R+�DI}l����g�򇹛�IU��Ʈ. m��XM��g���m|�!�����J��_�{z64EӐ^_��?c��i���P��D���O���;P�p>�hZ�g~1���Dd�-��v�Yζ�b���S��1sL+����E#e���S�#y�V���ܷ� ɩ*,�^��$�&%��9;?`���7�e���^�)����+�EE--;i6X����j�(@TE��������8�?Sn���U�^(�aY�f	f����\i9�=P8S�,���C�c���TX��A_ �:9���
�PT�oL|��N�-�_�i�ߙ�lF|��;���P@^)_�'���oR쳼t$1�5R׋��ǎ O{W h꒣���L�3���ݥ��(�k�\�?6 �� �;���\���汉B
V�wtMn���~d@�/�K��WV��`���Z[)��͉��-@R��g4A8��$v���#(��b�&�nZ���t8Gp~OU5���}��X&!��������f�+*�ݙ7IQ��--��,��]�)����,k��$�"b�VG~8� Z�~�b^�͕@Ik�aY�eۊ���v�$=���<�K�fC��,��Z
�w�j�6�?gl���$�W�\�[N)M�:�,M_1��5nd,etO����%���koG=A�ch���4Z.�K#:����Ʒ�zK��z�b�2��'��������7����z����	����`ۜ_�0E�M(��Wք�X��խ�n�)A�_L��v
�7<�8��"�bEb8��P��e����T��5m    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
/  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-#�,�(�M5�Vt�2b�`ak
ņ�W��m���d�-H���ۂ�h������p����o>2|�񋁃��AB����@���B���ՂD|�kF�`ƪ��.���ZkCU�� ;��Z<�mBXp����E;�lf&S]%N�{O^1�}�
���$�A���O��c���$����2<}�������f��`+�[����0�$ѓACQ�/�nnf7",@��&&��w�2LZ�����`~v����\}j=f5`Z���7pp�~���0h^���"���`����7�`&����gX������pq6V�o~����Ǻ3h)K����Y0�>�p��[��y�8�L��)J�2LZ������b�4����2��`z�I��~�DdQ�'���\�{�Vpp�@�%��Mx,��dAN�BxД��2�K�@#�C��u�����8AOM�/�Sk�������;0[\����F������}��ӗ�pu�~��*p~v3&�$�^��a�������AMA��ƽ�`���6C��)\>�en&!Y �n>b�u���o��GUA�}p���v�����!���'��(��x,�PE�mx,��t(�j��з  �n���    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  sIDATxڵ�	Lg��3{��[��(7�rk�խ� l�
4hk�iZ-j�@#I�Fۢ��ƻm�Ŧ�B9k�6�ԃ�@Ud�C�v��]f�ߌ��(�&u�Iv�y�������Q��u>�(��/K=
���$��0';�e1B��X�t�?o���7�ðH٘���Ve�f��WĪ�z�m���j�����c<�R/�67l��o�KQRv9�KW�UQQ�ƩS>�@E�`ҟ�>���h��Mi+��]���+����^s�	v]�(
�Hf�A��y'Jq��A3	׹��WMTz��7��� ^�Z�Mzr���D4��8�M4̃�����Hf+%�,��aS&���e\���KW��
4Yq#�DG�v%-�A��6R	L=�8�-�P���7��j��X{x{96M���je�[t
�Zڒ�r����:N�zc���Smml��܁ҋ՘5= ��H���lh�E{��mzx�8A,������������}! 0!A��l������كc'/ .Z�X,$�Z���,����?���;�(�8�_�RߧSj��,�bW+%��ysff� ��
&y:����f�(9�?n�%q��KE���,D���
NB�Ԛ>�Yr���0x_�vF��2���)���Nt�Pn)/*�;~7nj�t��Wɤ"�V,=0%��È0h��l���ހ�[Z4���e:��ɌzX���܎޾�-�-eWo#j�TA�-��eڍv��?��G��5vr��{�'I���N!�CLllc#�(\�>��3�a��?mCO�fގݽ�v��4��A+2�0�z�0 <!Yᨐu��rpcG���2[�L��@�v~��-,�gB�M�L.C��[�9�O����2���Nc5�����@?���� "��s����F#���������+
gF��du��\�d�-�K�Ý�F���#I�S�.��������EG�
�+H1�o*�o���/�����h�W�ɪ}�M}��?M'�����	'���m��:�E���DO�q��d���*c��^��m�t���)�1�#���1h��3�ɴ�#�'�_>9�X2|b����"s��� '{ƈ���������҄E�n�3$X!�^18[�D~e����>rE�Ī�
��E博�G�qّ�&��w��������$$�JH�"1Db���������I^�ɰ�ܽ�̽9#/�'��.�����cW�
]�J�����[�@�F�VM]�e��� U�[�ڗ�d�P��#^81���)�;��٢#;��Ƌ}��_�B�~%�_\R��׾��o�N:��.�L�\+��9;��|e�%���u��ۜ�,,�[�@��1���;�/w� Q��#_�������a��|�N����Z��    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  :IDATx�Ŗ[L�e����T �)Th�]W�:��S�5fq�1�8$&��KMv��x�Kv�yx3�lc�,�0`09����@�"P`L�oEJ�1�o�4}�{�����~)����{��,{L��n�� Km�$��Z�'v�$�2|>���*�?{
EE�����P_O��gc
	c�������K�:����:�Da���su�왮��0�L���w�]��V>>������K+�|w67[S7�"MP[+���2�|�*1~��L4�X4�?ca��=�ӝG���
���<,���
�=�'�����c��+w�\.�R�@ �T�x���4A8��}�׌Lsrw��d���q�����?�p�7��x>�ѝ�6���?��!�� �Z��T >�q�<(++����E|&��F�E ��lPJ��T�e�3A���cC��rYL&;�k}.�˭��A4�C�mN�abDw1��:�	��%�i�b1���JQۯ��am�$f��m�_$�<��ɢ7���gj�
�Q������oaq~��N�m~H��K�PJ���	?�y�|�@(�\(�]զշ��c:L�n�]�0]Ô��V+��fA�/��i�[�ֲ�fl	~�>�1�o�"�@Y�����6#���.�3=�Y��kd�
�f?�k0fv����P_������C�Ԧ̐&�~!����C�h@�T�@�
F��?��寒���ds,�]��'���Yܸ�5�ܞ�[,G�g��ݲ�2IJ4��dK�S�͡�R7y���i�vPk�Y�>���K�`Sր�^D���d2Χ���˺��G �ˡQA;&���y��_A��>N��|J0\\Q�)�8M#p��ϑ�;S|i�P-�k���A)�����W'�0\���h��I�_��J���ȳD�^���s�����5R-�F �B*�D�����\�yRqğ�/���76
8�H^~�.�s�����g�$��"�Ǻ��o���O9���TY.�(ؼ_}�b����Mcna	o��4���z�O�+��'�Aīږ���w�)�ѣL1��L扇��"0�'u�����C��B�R    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��ULSW>罶�@�ө��\�D7b�D�DZS)���1�$�ef33��e�$�L`@hujdd[�aa1��*��qD-h_�=;E���G�s/y}}��s�{��}�!<�5�b'!(��UX��X���m9�R�:�
u�Iמ�0 m�9������=΢	�n��ɏr$��T�HR"l%����:����� ���ǅ *�E�n �4��> ˾%0�k���m%���&gQ� ���t,�͜_A�s=N�ӏS�M��q�L����{ mp�
���j��Ik@	&��;�H��~����zݛ�`	!��� �V溓�7��
2�t�t�{ �r,E��xM���!�_����^Jβ/�$86������ �}�PM�����}���تI����������rr	s��_{9G������nO�mA��ֱ�.�V����j`�:�8�ɲ�v���N�\�e��ճ�t��e��Ge��b����*�r�ߢ$���"��㩊�c�ǭc�9\`�D����Y��H�O���Zy~ob=o��D���FKt�U��jVJL���˥���	���,��և]LQ�~���F�׃�{K*-�c�C�*�}�3/U�hb��<���OEEAȞ===���kӒ�����A���/�Y�zb�I֪�:9�BBBD� �����L�����\j^j!\�.�L��<�?Fs$y>9�"����Wt�VgyLL����X�1�N��}k�����:��^A��@��x5"�H���7U�5q�osx��L�n^��E�~7¼!�	��cu��%111i||h$b�l�9�v�,�	�����ƈ�l�� �Z�X��{��۷><�g�ؐ	��V1%�*E�ugf����8fhq-����
��;�åR�ۦ�<��(óZ�s+a�C^J���_�h9D��f�����?I9�m��[L&��}p��M��o)�YV{w$6�f3�9T��yvZSd��ޒ�v�,Kl��u?�}�i���������@ x�ju�un��:�]��W���7��e�y��Կ[�?�t��8��d�a��k�th�t���@uv��]�so�Sxj�	��[�7�����/�6T�zU�o�=<_YƋ�>�7���	^ ���'��2.���x*��Y�۰Ks'�}���<�JHE|�5�07�f�\�W9Aa�U��f�^��AnỊ"#�(aK��)�G��{}����h	pTN    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  VIDATx�ŕmL[U��脌2� s��Rڵ�uP�
2dS�,C�E�%h��Ĩ���c���Aݖt��A� ��ޖB�-
e����n%�24�'99�>�����9�r8�/�Z��pxd��quҴ<s��� ��򓈊�M����Bf9�SI4*ߚ�P��'�Ʒ^��l��8�������OP[�x|�u�
*j=�lnܨ�^�p��v��nחT���}\k�y�ˬ�5RĹ��:��&�<ׂ���!��Ñ�BL��'���&�����]��h4: ��)��n�/��(z���Ԭ�
/�@G+ls���� 6��^Wt&=� 5-	q��- �i#��kf0^���v���T*y� >���@,����U�^�h�� ]0��dŲ}��46�چ���I�Y�zӪ��4��X��S�7jr�t���� ��A��o� ڔ��llf%��,L�a��S�[�-Z*T*E��M�z�0��TM-�v0��ك_�Щd�Y=�n@SpXT���a?��[J-�&���ucB��,�Yhj<���.?,��@�!+������w�h`g�Qr��H�V���irC7����=��/��Ee�&��V�B*d��I&~�ri�����U ��
dlZb'I��"1
sR!S��K�yXuCv6�Z__��\PWW���˷�x<
GΩ�+- y��w(Ke�$�9ĭ���8�����L�S�TzFhT�l���,^��F�Yap|�	�����e2���z��+�/�ߦHW�~,8�#��,���ػr�0�;�E{.�OA�/ǵ�{3�x����L:�T:oم��%������E\QR��Pj� ��Pu� �6j��Mhu���'�Qq��q	I�yH��B�5<L�'�P� �RJ��Z=kw�OR�U֠`��ة�2�{ـq�_x�B���ѩ�D�jPRy�!�H���w���{��9(�q��!;#��ҽ�����p��C�J� �EJ�E��x�x
�[4(��p靀.2���u_�x�uU��gj������(�#���������W�Ƿ�5�W�?���vR�����{u���_��Q�aK��    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�c���?-#�-�%�ٻ�*6� �g����~���oO��͸-H���F�?����hcAZ���3K�-���$�[��t��M���w3�ga��/����0E�����*d���|L���������Í�W����s귟�+_���ڱ���� �/?��mA�W7/���2ܼq����Ǐ��cHw���mVe×&���8[���03320312�{�����|,_���00�0����u�031��3ܸq����G:�F�Ե D3��n߸°i]<I�=x�K�����͛7�?}�P���B�J��`Z���{���.2p1~d�����Ld�A��A���u�G�=��������k"�}��е�(iGX��������_���?��Z�ni̧��%�g�F1���l�����G����ϔ�xI <���-Z����o�-� Y�K2�v���u�`�V#��0+�}+�XP�����8�7���o9n����ւ��yԩц~�Ok X�xd
�)    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  [IDATxڵ�[lSuǿ����6Z�^�2��i&,1^y1t��`0�!����0uj��^����A�`�hI�!111�d��E�ѮWڭ�v����n�fg�_�����|N����+�q�� I���6��U^��>p\{Ջ�p{�w�H手>�+%�/Ɩ8v��b��wHj�Z}+ԔMr��g*e���e��K/�Y��@�[���Ň�Ϸq*��:`�vA�TՌ+�"��\��lV��b�6G+���ף��s�v���l�A�Ka$����ڙZ�������'b!�#�Q,�A� BZ8�񊩭s{��~��X �����O���Q�Y.`�� f��a���L^}�8���!��t��^8�1�~���[.�CWZ���OCO������_��d����7PH'F|g^���<F�Ŏ�'uB~פ\�c��V5�	ǽ)ĳ^�p�y�h���-���|*�o��E���v�D@�gH�k�l�Z��}��g��L.ᪿzI��fw����w.�o~-����A.���;'D�c��5[����7��t2�<ІP�ơS�ˑ�$�B|��rSeq�d�_.�@<���;�)�ܰ8�}0=RR�g�fC8;�,z�:�J,�>A,M��	i
��ݼ;�|���<Y{w��$Ɇ�Jr?}�X��
��&��_,��cY���9߄SWغ�hn���رm3�GNGp3R�� �������{z׺SJ4J�F��`�|��e7���Q�z EÞ�[L֝Bw6�~��<;��L�ڮ�J�C��E~�zM�t��M��)2pK��"ɴ�f��$�ar����]�j��i�����4��NW�'.����3��d�
?�|y"��j�&���!��*�����Mұ�������Ϧ��tUr �Eq%7�p}.9�t���ְ�Q!#qlO�X��s�H��u6�lZ���N���R���;�]
�H
�����.��g�Ǻw�&#I7?�(�MM�������T*�h�u���
��6\�����h>�8�T�5
��_�r�d��gYF��+W�|��J*�u�{�n�mX�ե��$�A��G��^U�y��,�y��?�Х�(��bU�Y��    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
h  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڵ�{LSW��mhl�&s���b�2��0u�d35N	1A� n��m��!�ԉaPж�k�9$�nc,ۜn�&+�1�	�(������SRJ8����9��|?��@���?�v���j�;�X�O����9	�4y%�)ʳ������mp��[��#Q
��-]v���g�H�%�w��4dǠu�m�d�U��n  �Z~�튄�%�����yZIC[w�պ�<mC?��p��Y�38 L���Ȁ�"�.#�Pq��u?���������(z��c�b
�VΆ@�z�p�������ؾ�4C���ȉ}�`��-��q����!�D�Bd�1m&ּ��*5�ͭ8|g��\�D�~��4��h�'�ކ��f�+��C[��
9�L{���ʩJHr�ͺ5�ڝ(��4��-���R�08�Fm�e\����x��l��Ԅ������@���lc{r��O����}Z4(p�g5�#*�p-ܒ�`j�U�W�4z��Z��G���_C�F�[]O�/�}�?Y rq�]�yyY[�-���o�;?�!��������w��G,d
��"�E��&�'O��b��;G��!sS@ ������b�@�ǗHY�f�Y\�Ѳ���vH��]"�$7A��5���!�W�,wH�TC�V�7G�P<��+��~h�'k�y~Hȿ@�@�"��/+_�fYBȤSU\���Vy�ը���m9�!'�[���k�X{�[4�Rľ��+O-awms�M��]��.���2�~�����@\�9���NZA�
��E&���� ɯ*A��$����Д\D��|`k���Kd@B�
��G1�~�껥�ﬣ?Q@�3o`[D��Z<�em�8�.ؒq��r��G��=�s�|ka�u�?#'fM{a�܋��V�R����c��# �$���C�x��    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  )IDATxڵ�kLSw��}��G��h��a4�a�Y�,ӵ�nY����e_撙}X�@��ٖ�����[4)I�Hbܦ��(:�!ho[A*H[���{�ν`yL2�|���������9�s��$I�,�X���ڻ��ʦj�Y��<���O�����$�w�OH` 4�9)I�5%�~iY��a�j�"�~��\76�}e N�5�CF�JJ���*�i
��D�a��}�L$.�9ʻ��͝���+�$I����|�����J���U��M�j���B'�MOa|l4.��o�z��M-{ ������y����6�'?O��4s���vy���#�Ǣ�\WT:]�2ha!
��1hx�(��Ѓ)�7���V� �y���Pql��]�G`|tC����/c�i�;��+��YA�Ѯ9Y42�wn^�]ֶ@���rR���mch�V<�{+.
�7y��Ǖ-��jg�q��N6�~	XF�XL&��k>��Z�����/-���oye����x�|��]$�l�+�q�w��������F�j5`�\�x�X_��|��;�Q��!0;�O芎��hްv���KTx=���l~����8��ٙ�q��W�rξ�X��\]�%���� ���3�+98�/5����CϽ�����}g�> h7SͰ ;�|1���g��a��3־��y�2z�!�0����i]�%TT6U1�ڈ�b�h�p+�U�Dsa�b��	gi-�h�f����w۾�-Ț$�jh�t����Lp��u�K|* ���
�Kʌ�<t�+���=֯�
���s���3TryZ6���i�$���n�7[�w��p�Ui>+җ+kB��!�f�r�8ɧ��=��� �vpƖu^A�6����J� �N%�A�q	��h�g"��S߿�� E�Z5�3��}�.�Ze]AȂ(8�f2�_���7��k�V��n ��X����i���E )	��-�i���;��Ɛ|��70�IR �X���˧H/&"�T�l��<�$��6��~Ey�	b'.U`�����#��6��=+�ݎ!�Uuf�    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATxڝ�ILQ��#X#��U���z���(P�ҍV1��rr�q=�^��h��h�P���
j � v_��g��N�O^�7�˼ߛ�_�$70�&��_j�U�����F��N�o>|���`�t�Hu�k��uvF:٠UՆi��?QS8� @.W�Auf�np>vTj9V\�Z�´5 ��@�݉�{B8�9H�hԁ2Y�6��������١	�H� ;�wq��� ]�60@,��l��J!w��
��i1c��䋥0Y츼��콨÷I=g�츀��'��h��HF�颃�Vx�
���´竰�II� 'O�\����mX�
777Q�0W��:�G�a�*���9b�1R�����d�+ZW��T*ZaU�s
��1c��f��(R�/��ϱ��eA+ܮn���l�����2R�*�11>kX�
w���%5]�3Z蟡��j���&��"O$�Wa9�H��N�&���4liĭ�5����e����sC��c���p� �����Ow�(��S�=qC��f�<�Z��d%B��\����NM�&�*491�&d��0��u��"��wD :��k��dƻ1=*O#��]���d���Vx�0?.���a0Z�a&���o��d�W�)ȟ��VV��U��9�#�wo�g�чz��d�e� �%��Ӷ��Z�Q8�U8fe��c���A�묤��p�? �T�Py-~��SY�ݩ=����d���X�����~@���0s	�)�P�~��m��޿�Kߙ�Ї    IEND�B`�  Left(Top� Bitmap
      TPngImageListEditorImages192Height Width 	PngImages
BackgroundclWindowName	Save filePngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  mIDATx���kHA ��z�'JP����`!(ie�Q�����;��
*���,�Ea��iP��0*(ɷ���i*�Շ)��y�mo�v�ֳc�/α�����ff�;� X˂����@�j&$���Z��\�5���j4`s��~����+US��&��J��8~l��Dy<����
�J��?�J
��X�=�F&vJJ&c�4�����1��'��Ԛ55�h�Z���F�r�/,l\W[�����l�R��:t��h@J
�P$��K+7�$'���LO(��hj�CT�T0��#+: ��qW��T�(�)�`�'
��з�Ѐ$e2��	wӅ\z��[� E��&�;�[ν��e ��d�[0S�4aN ��;���F4 A��Y�V��
��ф��U03o��'�D��[A*���'���+��jF��J��3	��Jw��ìq� =�h�,~u��� b�`j����������D>fG��b|7A�n
�Byk�ѣѱ��g�2s����. ���%b�Hp���o���64@*K����I����d ��l��F	�v��adr$���U��[��@;%S������&!-T�]ga{X4�_�d`w����Nl߽;�H��ǎeʇ�4 2F��IU��cޓ����R�??~�곯��.���nv,SF�u���]e�<Y��r�ҋ^����FPwN=�޿��7��˔�C ���m@`H��Ë7��q�؏�Y4/�#����o�2�W�|�.�l����������rs�]��lb	 w
;N�V�0�?#�0�_0�S*?��vX��;%kQ����=Ib�    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
R  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�ŗyPW�B��Xƀ�����E
Q�:X�j��4v
:H�*�h��2#=�r�::��%��B���"8j���&l�����"���'�{��}���vCp�A��*��s�G��T�-#���g���� _D�WEʦ��,9%�v�8@���ks�gD��� �9xPUV�d�y �ju�����h�K��)g<"�����m���p�zgl�,b�'�=�£�)^C��"8w���� ��AP�U���|��2^�B
�'�b��!F���&ڭ4/��1 r��5�|�F{`Ƽ$O>�_� r���I�`W�a(�8�U�-C��$T7���$�^�:`nL�x��|��3�������׍f�w�8`�j�dİ� ���]]�m�q�~o�t5��e�#m2��[����9��UI��Ç��V����W$- e�37@aQ�O�[R�����CRW.�xy�AT�*�:)�3���{P][e�~7͌�<?��Y;�$�Ε�);����c������O=?U��b�~U�-�XW�W�&��4�O��} Pi��$��&�c��} ��_�#'N��s��f��^�}���$_��G:s�p2g���po����1ӗ8 M(�P(�Аq���q�q�N�C�8��h��E���wP�8A@���ӧ��z�� ���o�#���:8-9~��
f�Z[hn~��+P��)t/$~���*�=i�E�՚�{yd��j�O�Թ�_�BZ��ל�G���aS��>�&��R�:��s�)]���7A�<������pQ�D�k���$���C`�oep��5 �A�H����`�ouELg�P>)��8zJ�W+�U��Tr�>�{����r̌q���li�k�W�3FY���,7�X�)�jDJ���ݽ3��y���c�X>'X~䰀0���hj�
u'Q���Pj`���d�@�<��-̈�7@��url'�J��7�9�e&�_�Td� x�A푭clًrL�ihVg��R����e0�c��T��gۜpt�P'>?t>��X+Sd��<�����ݹMw/+(]��I8k�2ߡ/rimv�] d�2 s�
��<h�̑O��ɘ��<� �ޣU�����5��/^,&w8���C�.��Q�:q�H�۾ނ��f�u-��=�\^  �_���(�&�sؒ��T�e���9���W��S6� x|'��jI�u�5Ϯ��I��j�bZ���� �"�"��=*�����:{@���r�cѺ��o Ks����������Y�(]��7����m�bi��u/Z������4��[�Rt�?#����OQL@�@L��Q1=���Qu�q( �-t!E}�h�����Q[)�Ō���ˎ�!'��tT�����=�CMvSw��x[�_'-�`��    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�ŕ�OQ�O7�����q�QB���>���n4
h��C5B�
��"��QQ	$�� 5<
�o�-ס!���tF��������L�W	!��6��G��$!�d5���J�����w Jt/I��3�S��#�C��:7o05Y*����r�,"�����'�ѩ�c˾PjoT��/���9�G�|�sa��k5���_H �f�*\����'���7`x>�:���1x�!,��� �x?13m*��"�j�3�@�O�WS�1�y����>�
���� �NbVe�����D��{��a�}!���Ck�%� W��\!�'�u�v6��3��0;��Z�) ��N,U2���>�(N?[��h�ȅ��� V�W<~4�}J�!��� 9�.bQ+��gp�PG�#xע+,*@��)�h���O܀�Os�(�
�
���` �����>La��=
��2V�]q ��6b������o ��
�ٟ�PY�I���:�]�ԁ�hA���
�ٿs[v ��b��a����U���-�
ˢʈ�����:�Lf������+��J)@�a�7`vA���j�I�����g\�bK����1�� 0t����HO��2�Z%�Ϡ�KXlQ5��I��x �����U�¢�Dvr@׍��� �
+���R����.O8����SX�+O�Vu���|� ��.a�E��D��� ��&Na�R(;[����P ���r�� �֞p	k���+T���_6��/�.    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���mLw��i�������e��_lo����(�-PQ�2���	�([u��DEJ��V��d/��D�\a(���B��Z�+��9�Q������_�\z�=|򻻦ex�G0��T����`�K�I�����������L>�2�s�� Ti���A���cC����L�?@2�������~�x�ؒW
P��]N>S��"�� �+�T�$�~RUL��J:_
P���:���D�d5��5�LBSvmO�,�>�~���=4�8���k�V <[�v+�,�Ȯ陱ZI����#��B��[p�D/ �_��鹾��G� ��@������OS�O�~�|�Ƚ�T�v�|�V��GxXL�p��(<SJM^տ���f��	�� �HR�f�'	0.�
�sc������ �qM�=7F���&���%)a��e������1�`a��ZK�_<�ޤ/�j|���Ho���I��<%<\ e�nIώ� �.��'��e1�� x���`�؋�|X�v���]���󝎱�zF�����$�_��I��3�ӍͲSd��E1�D�}+*4��OTq� x�{`8�Ƹ�/kx0d���Å�p�Z�2��v	�� rP�m2�����$��tp� ������6j�u��	 c,7�#Og¹�q�ڸX�3K�)u����Zᘯ3�R����A��P�lT���
o��zT}�]�&&��^��	`lN����'y�c��<��OD@_�j� Ȃ�(#�m���5?dP �Ѱ���>���rm:�'|(��"{pζ±����wR QQx`PdB����xx(�U���]�՛7���B-�|� (+ډ!�C�ϲg&��Z�;�)X5�s��8�U���B��0����7�^�	��Z���\�,���9,�IN}���K48A ����o�-y��~�H�(���ef��o:    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
5  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�͗}LSW��}�B[Z>:�@? �aE�2]�%�8-_ۄ��%�k����2�lY�gm��k	��Kfb�	�b��Q:����*��k�Nҩ��L�nrs߽����;�sn	���"�� B�1��#����r��N)}��7 h�&3C3��IG[͵��62�+�$ᡔ'P�'�a�P�o$LZ�m��m 4RZcY�|%5�߷���շ�7k�&#�Ujj�:3K��TH�H!
�Ϸ��ρ���]����\uw� ٵ������������dÇI���Ţ�\q�pw1������r����*
`m1�o	@��yX�H������v�3�w��xd5G��;/�0ꪨ�M@"��XBT��t cw�R�٥�S��[�Prr��	�8��y`q��Z&22U���z��Y���~�M{[��M��rs��y����3���D�タ��+h7
� <N�t�VW@�r�^x0s���_��[��3�.�
�fd���-���a�����9g{�Г{���HK�J]��/��ir�/���ks�相��k���-EjzL�������Ϟ�5�\�g���ڔ"Fғ�K�G���� ��y�?��w�����%�,n�-/-e`�_��X3BS�Q̈$å�����Q� ����6U_�	�.�/)?�B�̦1�0?�1�L�8��ۧk辢)(~;U�)�g=p�'��6>� �Q�)�I�J���4�\��	�֟bZWZZf�:_/�}ˋ092pk���� ��ɒ�]{*b*c�~Y�0��#�՘�c���'I&�Js.�Qs�g��j�����$ٍTen�}M!*�1�|NL�.���>O�]C������4vgȘ����������  �Z�ɔ�[�� ������ao��ߒoi�'/I�i��5���񡛱�L�ϣ��?�OL����=tA lc�vtA4K�(���}^�P~�J'�WW��c�j>}�? h�tƽ���}b�TX���ޗ֖ӟ�8@��$%I/��}�M���l9���P��>%�:�*��f֒�[����>[��b�+ٿj�	�D��0�iل%��~��7쭆� ��E�L�g�h|,N��i@Qt���/Z`�V�:ж "7fJ��T�CXIR��T9J��%��M���+�*�S���*#w�m`��Hu!�S����.��G��Z���?�9�Qw����o�
�m��GѢ;R�"ξ��0m������K�����4�:����߸J�u��"u�S{��9��g��F1�HB�DDQTT@��|ǐ�qr���\h���c���V���A�_�<��b���	G��Q/���m-�Ӱ��E��7Ĵ��:H    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  bIDATx��W�Sg������d�E.!h�:���k�Ҏ�N����A}�S_�N�؎�δ�K�A�T[B�Z��H�*�dw�^�}��l������~����~��a����)� �a��x��"E}� p5
^}>���0�� P?V�|d�wH��K��ʫ|�����G�����o�c�?��Ł�r/x4feAl��3�@�yE�_I�������(�ҙ�����8���;(�5�..m�V(��D<~0�6
2 �7�K;/����Uj�6ן��FXUQ�G{���<Hqi���[��!/�G�A"�ry8t�K������]��C���c ��A\�S�����r^�tƃ�;e��<О���>���>6�����` p��� �ˇ��`�<�Va��ǖ����9U�"C�f�9�Y�Qq^a!St@�?����Ź�\�=711�ܑ�u͝p��r��{��f78�-/���脒d���@L��DK���Su�������Ks`iaz����{}k���Uu��m8Nܨ���8 Vg��0�N�h�io��S���fwh���-�N�b�Zw/e�9d��p�}4Y�
��~.>�aa<]8I�੪����?�50?=�*	�ɿ��֟�@�>i��+.��9\E�械B�aț:x�ɜ�}C�;?3�.�R����&����tj�	��]Xv�UXb0��8���hM�s,L�$�����`�.�"{�Q�wc6k��Yx6�K��X��%I���=� 	j���g+p4��ʲ�+I"���*��#��+��� �w�;�N�����s�����aڿ��kf������%;f ֻ*+���&�9��,=V�����LH�yHJgx(x��*�	�7[������Ρ�A��1[b��U�aK�(�>��Ua��2P<��]��Ŕ`$Ei�R[<H���Il}�>�AcgIb�0j�0��$7�g7a'l31��H��T�rS�~��s(C�px��>�rς�v? �v��J����	�M2��X�~��Ϙ(��
vs=��l�~x嚆����owR���S�%7'����Ӱ���	#�^[��J�@�<���߉-��ɟ=;8��y`�H*LO*�\B
:�ȹԶt�1�v���資ڳ���Uإ�H$�e 7"���d���i�����J/5-m�I@�2��<����!�ǧ?ͺ�5���Q�٫�GY��]&YE�ZG���9^�Qn2㽐�>=�	I/��_g��˺��ɋ8 �x��9Qj��`O�^�k���J��)�6k��R|"<pә�2� ��W�$U������q�����m�N�dA�GpL+;�4��͖�.��v�l���/#��G���S9����m�� �i�
�3���    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  rIDATx���{PLQ�o�^[D�d*=��#�h��c�ь�fL驄J�0���˫H��P�͘A�`H�I[
���d%=��������=�=�?~�����9�{ν�h����_���"�g�ٿ��9�1&�bb�Z'��9����V�֘�܀����� 29 �}b���m+�;����Y����0�l;�iX��^�+��C�5B�^)@�x��	y���񀽍�j�
 C@�كؔ[��2��h#9���i��	$ �j*���&�ϱ���!��Q��
�����:7���c�R �Y%�L�����ɅnZ+�-��W�����-Y8~�n 86�p�` �iH:ys{'�?���+֯X@�d�)���:����!��D]H�o �B��u�6�VB�*b���e���}�P�؆���h� h��g4��LG��j"�-�83�U��
��FzSWfޜۼ�ȇ� iq$���	��
�˭�<�Y��KO�B&����܉���T@ ���3�{4W�;S&����=�f[��P_���_����J��* �܀�J���d�~̴x����}��.�n)��Ǵ" H`;p*��v�Ee�L����[��tO�m,@�	O� R� 7��QXZôyz:H�����ӂ���PK�=��=�*� �F���Ŭ���1V�9A[k�_7�Ie=�eؘ� �-	8D�(�$ĝ��.�[�:�Z��Jv%��!�v� '����'\��|֗�榓�q���X5{C<1�ĈU��p7��
�,dw@�ӗ�{'��^�;0m�D,r����LhH�|PR�
������]P�* F5�OED"p\̀H��>���( ���#��������H��    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
Q  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��W	TU���܉;1�C׊��!&����F���ӕ/�x�zM�d)���e�e��S3�� �J%@@/ w�^�|���o�H�V���:����o��8�̍!��U�bE��ůܯ�Ҁ�>�|G�w����M���������p��u�M��pk~yI~�C S�͇�kc��X���_ʫ�(ɟ���HK�#U��8��zOqA��ټ��'�|a���{���p8@"v�'W�5��\ԧ;����r������2�m	�p��G�f&M���u�:zz�����8�yub���	p_D8�!��DG�O���Z���;���1-�e�H��5�m��-m��폺����LUqZ�L�c)��d��H(��������ғA*��dà	�8��2 ˲4�Z�a��c���3�ŁP$��������"����	(UU�֭�����z|�K�;z� �����t���ڝ�Ğ��_�&!"秚�¡�ՕH`ڨ�fG+}�-xs�k���]���Z���.^RSB�:��K@8B~�n�	�`���v�M���T��1Oe�����X�E@�c�����w@���N�a88����:��A���C�׽���Jhj��WQ�Ϊ1eA�2{����]�>��^/�����YS"��c����r`���b��1,����®�ЭV?��dc�`�9W��k������`�h�9	�� �2���l�3�Zqwu{O���Q�|��B�5�V8SQ�q[)�+"'��5��Y��:4����UBf�L�r>���~~:�B�ܭ����<=䔈IX1C(`�3䃒]p�O�Z'�	�]�2�ϲi���2���)�'�, qc*EM�+���w����-�c'1$d�,�D���I�\F��cy� �OH������z3^�0S�$�>��N%0?+G�v�RwE�/�d�[�n�������oF��d ��a{�~h���*T����	w�9g�4�v��R����a/�z������p��	��</J 5+�����c����<߼�sP�>,�����u�@o��(~�ە@r��$�Υ�3�B�ぷ�t�!|�o��sk�1�ae[si�[,�گ+|[�X�O�.^���m�&�������L :��<�y%�:��/v���OwwZ|tz#X�x�X=�y��"�j$��Ϸ��ju���)�̢ n�_OP����D�������8�+/���U,�4�8��Q�H�#�Kd1�N�k���|��{��C���V�����l�"�x���O,H�x{Q0oO9�D���^���fUc��:��q�p'GL� �ղL��4��/t¤� �h��޾~����::�7�����w\�b��.���
r��-�ۣ9o*D��˗d�x{y��rK,���	����Sg|����}�Mu���k������O�����T	�#f�W�X��2������eo	NV�"� .u�a�f����m��K��^��)W��7yb������F�gR^� MI6>��X�[��n�h��	N��(��g6`+~��%�I�f=ΐa�	�$"�@.�;�3�,����@�����N��Z�f��0�w[�� Ir���{'��>��G*2��C�<����>�su0ct8���+�ΙA]M���'jii� 瀀Q��pt���J��Ғg���
6�Bé�숙�p�!�I�!
?ə��X#�d�G�	�� ���hU-4�؄ݳ��c\�L*y6}~"S�xO5�m(u!��c�R�ݾ�εN�X~�+��܄���s��6��=�u�OY���5'�ֳ���i,�F~L�2Rc��C�@��x�����1�-�5K�5U�Cup��I����kF\˰�ΟSԪ��٧���?s����Ph�
    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  *IDATx��{LSw�����U�����B{i-P�`|�l�",�)�=��h�͙���N�%f�e�,����=t>p[f@�m���	H��A��n_0�~� [�
.1����ro����s�9�sZ,
�bX��8рa�i�����Y�)�C���?�g'L���^�� �,�^[�*u�&r@$�ڮv@f�tii٩qIL��'�A$���؆��d4Bscݰ�Ԧ�p_ ��}���qp���pQ��w��Gv�ҕo�%+Y����׫����E�S`u���.�j�[2/@�����`B��=��|p���`�tAF $�x))L�}��H� �̓�����[n�|���~?(�J�m� q�����in���$�P���d�ȘF�k�n�Q�:[�&R�B_y' ](Q�$s��U<�� �F�p�Z#'(�U��G d
�Oe�E'V�U�	��憳��7��� *@wG�)�aˠ�>��K�r��������A'�V�!9�	��\��##���� ��6�\��(�G p����붋� ���a�|b2h�FF@H\Wo�(N�	h
L�>��ɟ�zm�L W�杉�l�=���A]�w�݀b�cm�$�9���2� 4Z3�!"S�K�1+\�F�:�@1�C'z��p���~B��2 C(^ϊa\�r����O�!�F.�V0�On�a��2�1W(y����z9 (�赽3R �a�'��}
�Dp���C��z���	�o��A��\ ���p2��vAIyT�W/��؊ ��LA-'�_�T��2_2qhLHlh��{��t~���KQ"P��Vʋ�F��ܼ&C�phf.ge��K�%H,�A��@G��b��-���[��ҹ P/щ�"�LՃN����$*ª���K�֤d
P�	����`���{�b��W�(�Yߎ���+^��9���t4����Z�4 ���d�$�K�#�ybH簁DB�y�^
�~�ģ{�wrG�FKD�qq��F�R��>�~���mE&pĦXf\��ʁ��X�� $�E!q���M��v����ňD����tB�jh>��Ku�#2��`�������c�z�@);�ơ��A?�#���f���ȾO"�/ �g���)+\3�G'�l�*T�'�����ß����qP��������x�8t=���8����H������U�zh��*�CFRs �ڂ�BBQB�,y��ƀ�f�u��)1z�����x��� ��
dK��0�y�{���:	 $<y�u�t�a��e��b˰M9O�����qA�ųz����gf2�0��Ue������gB�zMd��WU��N�k��r�/�>�t�u�B�R喎1��1�@���p�>��zO*��eS�RC>!���'#��v����B��^�~����iض������B{,�I����J!�M�
�}�4w�NjѢU��+����
���[ç�:��� t
f�}�Sh;}�h�������;u��l��/6�� Q���cw�    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
'  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  ~IDATx��V}pT�?���d���� ��%YBj���X�D���k˴&Ѷ�ɮ:-~�:���j����$�)f�°�P�&���I@4JB �~�o߻��B6�0-3��ofg�ǹ���9�s�a�_��N7�ߠ��ɾ޳�� ���,s-b=�BHN'NAN�0�m���m �����K�Sa�_tz{�@������
h�e��Q��� ���[�b�V/Be&6�sF�8�Uu]QhQg����J�g�f04�rbAW�� s��/0�GX<����I@�Z<Jevy>��{�@�������~�#���sb�>�ӓ�<\��&HP�������v�XdEY��R��uq`�����=銈1q+6
����uyx�p=�{�s���WW�/�>�=����O]�
Ŏ����8�F�Ր$ˏ��^���l�5���C��*������J��������X^��):�ĸ;���z{{Y� �`7Br�Up������ r+�	{n���vߊ�&h�Q$�ޮ��gǸ��qP`��c9P�$D��O���/L `+�M!3�al����M���w# � 	X�o��0����;�N<0>���9#0���T�W�{Z�#��r�&����Zǈ=����I���^���	�������#G��5��� (~�X8�����>�yjKRbn��o*Z�.u�>�M����G�e��E���"#'��];<'.{��n>��[X( �E�� �T��M
 �қHIIeHI	e�͎vu���f�ȄuE	����� rKT�_4��0_������
N��=$+[Q?��"F��]q��9��9CW��������^�b���6;��̩�n�	�j)*�?�my݀��z�����D��C���|��9�nڪ|>��P�D^��7���)b�NO�X���P'"�MJ�^�����|:v��s�͎�@%�%�2/�` �^G�P���bh ���:c����,:��1����O�����-N P����h�e旦� t�D���������=Gg���o�smq�{� �'�P}�����@�I�+M����c�$h0�ʐ5�����N����,z���ˮ�f�1�����fcZ �4�z �]�G.��Ct��ԇ�5(�1No�*1��H��H�Z<8�G�כ�?FuY��bj��d���w�eZ!A\)�)��֙���׼0�a �N�ή}t�����2�/����mĐ}��.�6(�peh77�F�p �	Y){4�·�t����9)?}�*}/�i�Ͳ� "�� B������B}�,���xt&dD���S��M�jk��`6k�\5R�6Y�cI+��	{ۓ��5B^���K
�g_q����_�������˒�;W�	Jj1	��gY�B6�0�`1�y��f���St��
�i��jJ7�O�:g�4�Ŭ��EF|N�}v��_����UN��M �����@mL�&bj�k�f��@��:5s�uF��T�/��v���x<�kvbO-H��v��8~�BW��xt���
 �)�8 @\3.3&`��6�:݃xza�/�"�<#){h�r�e��ה� ���_��w����q�"�Ӆ֛�z�4<�K�\����!+P��F�n4$�����哾Z�~
�?��<�O%�-t>l�Sʙ��[LͨXpW�BucH��~�(
U/^sSj/w=Bk@��B��͑��Jݦ)����R��g����?�tQmF.p&�k1�c*g,�Vx��]u� ������ᅛ �]�����yv��J`]-J�pk���~�f�dz���Q lC�b�gf�|�@ ���򒥮�����|P�N�/��<R�Fi��+ݠ۟;Z<�#g,�%(��`�N 1�Ԅ*�k�3�O��oJ�Fԝ    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
F  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��{lS�ǿ7	!NH�!/pb_'���&BHiiyt�TT-i�h٦��i+�[U�ڪjj˺V��?m��*�vQ&!�<JL����w��c�&x�ޖ4�cZ����~W7�s~���9��3�N���|/+X�_�0ߝ��`���ZzL���D��Ā�8��v���{�`nMS{麶v��D0��0����b2:Y�v=s���Ύ}���Q�n�`Nw�3������޺���0�9��c���b8v��=��Ν|oh��s����:���$��!�
�]��~q`q 	���a�=Xdt�{~��G�?���y �B�����U�PWW ;;}:#�~&�aĢ!�0j5���=۠�W�sz1����UF�P%���Y�X�/������E��B_�Y'�+��� (gYvY�
�'�Fi��0�%b�]fõ��R���eg~|�� ����ES̏�^{A���W	����� ���_-�9����H�*��QV�+�QQ���������رuӂ Ƒ��]����W2dʷkZ�QSz$��4��|��:2 �>nlۼ�������3�&���3�*}��]�ⲊE�0	c�84-H� �J�!.^��=v��Q:��YP�b<qW�"�π��h�1I��ɷ��}Ә����jE�(�T�I��28��BH%HN&���2*x�X%�y� 7�BE�z�$Ɉ�"�q���m(W���l��-h4�]S���1�lN�c�'�0Q[M#�qX/��wR���GZ6~s�C��:��r��d�ʃ�e��6�6�aM�zG�.�1A氙02��e`ޣ�B>R\^�_���1,�C0�|�.g��hvvJd��͏�s-�U�8a��y�8}�|�^>k���@Yu��Zm)�L6U�F4�e��Jjx��.52u�U�PԷ�Q7���N��b�.��\D��d��N`**p8s��U�j��WT�48ͱ��4�0��|Y�</��(�` W��#H�(�	�C�4Ѹa�i���5���is��CE�d|��z�� 4;��}37/��\��[hoܰ��|l�`�������!b~�����ʹ��ƃ��1� PN��tiލ���C"U��^AJW+m�[4J �8�t�]�9�{9��/闩6/������e@v�,2�Ǎ��(��} ��n�[�� �aw~�����w����
��9ǿ��S
��	��zs�uΪQ��8]B1�zg���[)\�ǪC����k{A ��?$.]uP��QH*Yh�,
D o�H�  /���WNS�`�O�m},c�;���Y�c�rѽ���t!�kk2�+�D�~RE(�Q�(e-ͅ���G8� e!����O�N�_ ~N�R�� �pt1$�ô�����TZ) ,�� }�"�����B�٣B'�n�}��������ؓ_PTr�ZN-���^!�����PV��.�2��}/���h��Ʈmm�0��Q����Q�)� Ii"�W�~z�0lc������`�m�Z�"���}g��KA������0�ۀ���Ҋ�OlY�S'洡��P�����u�{�_ı�ߜ�L��N�Sl��47:;�3 ��4�����Bt��fP�D�,�!��R�u�Cx)��өT��Y[�� 1�� ���.��]����:z���� ���Hv���    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  /IDATx���ILQ����!��Oz�K�xP����$�H<�R�
"�
R0�A��Adioċ�$Җ���bi)�y�P�I���̻����e�7�B����������x{QM�`s�2�#p���T�a��W��e�P�	w�JY�W��x�L  �XOԩ�p��PԽt+qa��P��,X��}��B���U�Ui!sP��a�����ڰ���uu�K+� �e��J1�!��=��a���8ʗ������ϓ��Mz(��,���mA~��:@�G�.�ـ�`Y'L�!LNN�	�x�V������6��+�Guf��Ӄwcn���a��3���Eָ;�D��E��T��Y�<�˲0��0�Gg�N6!�ש_8��o|�Vb���P�C�V ���ǹ���{�o�ϋ�{�'�
��:P#��;�	wF|�� C�s~� Tx���=���X0lDWG�[���N��Q�}i{ F�	Sf��Gp�R�Tm�͹�w��jŻ�>�%V�
�g��.@+�rě��02b��n�9lk����ž���o�J�)>��D��9088 ۢ�_�ğ1yZ�YЊt���I8l2`rb|�%䪥)������&R���<M@�3��E����'�^��,;+������F��� 'JZ���%�d�Z8����k�a}q&�5E�n�H�l E�6z���¾$9�D�-�(}���h���'D�-]�Z{�,�2�#N��Y��h�#�� �
�T ��#�$kݐ&@[pE @^�O�^��������4�D���� ��    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
f  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��W{lSe�ݶ����-k�V�u/a�0�s8#QE�t@ܘ� M4D1�Q�0B�G�(��Wd�mD�Jf4LyL�<�W�uݣ+��z�^��*��Z�<I���~��w���9�q$Q� E%ܜ]}�q�@���K9P8-�Nx�	{��Q�����c71�=���6���|�B��\	F"�H�w�|^����vLڭ���z��}��ί�|���6e3b�X&_���B�P%�Vפs�ݮ��[�w� �_j.�h�5]�����	o�� 'u#��C(A��
F,�� ��-f��{�T ��������:����]H�R��'1:���T��e)*��@3�;kn��ƛl��{�nq�n������´H㼲���Ȝ%Ay�J�RX�tܲ�t�ܬ ��"�h&L��w�Jy���
� H��,>���Y�Jˈ����%��2;*�F���ś���!
�̜�ov�Ƈ��uWJ�Č	�PӲY,���(*�|b�)
`���;k�ql� �f���
�k��C������L=W�q;�4��E< ]:Â�<5�t�ώ��,��:��@�o� /e�[��%y���3�F���>��7������a U-�b��=+��hE��W��>��GF�#�������a�4�[b�1�^ô˽�����0 9/��Wkt;T�̘���d��2���6��:} �������� �݇�C�1��`�0֖�	�=S?�T"KA<ZQ(�\,�7�8/�!WR#Z��A�]���|�f���� F�/�խy,@M�PV~�N$��,Y����@��d�%��^�m_����nr~ˇa���<=���E�$zR������ao9�)�;o$�ߨ5c��Qv�� @�_�4 i<����}��\5y��qN�?��`��1 ��+��DIX4���-�A~���0�$���}��ܚ��5:�2�D��犕xwMP�G�/����������OU�ޡP�%�h�N�/������>��lRr�V8lc�א/D�TҮ��$��/�R�>g��Y�������Se��@Q{������y����X�8�?��BB㓓���5	e�~{t�HR~T)�{Avu�b�s"��W��b㓡S��>����2��Ax=S�ߎ5�U�4ő�@$��2˴! 7x�����L�[:�u��m�<emh*RL�Z���{Ċ$�X�m�B"ġ�16?	y���Gl~����~?=�<�j��"��w��t2]I�v&�+��>��Y߳�/����x(�nYA	��)�j�T��/�S�I86��4T�p����r���|�&�f����f����|^�~���*z"���Ä$�&��&�2�˂'_�apG �']��%.w��
˿�����z�D�**#VWQ�J�$�����z8p爺�W~�g8.�E�_�i�ߥh'�    IEND�B`� 
BackgroundclWindowNameReload file PngImage.Data
_  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���	P�U��.0P���LJSe��X�6j�v����"�r,��ASr.)%(r�G�1c����!r����뱋���_6'��������}��޾��!x�����'�[�/"��v��?1ٗ��͎7��b�������V*����#�P�ؚ���+��f�Ĵ 2�n��o��{@��!)��-c�H�����-�A�hC��]�V _^	߹b�B'�P$A-�FJP�o�
ּ��;�
H��[�`4��,<�?���TM�Z0>��B"w�@(�P{�W~��!�l��^h^#�'�'�g-b��nu�QTw�uʅ�m<�s_���6�mh���y�~e^p4W�W�o�����D����/���a�(m(��[�=}�������x�y'�]sG��Y������\�s���e쉺@b|֡wP(o�
�|m� ,�pQM�ш��/��TnNCb)�$��e��'���AϠ�����pJ���y+��j^z��Y��w�,�ץ��Zp"�5_�7�w4/3���<�]B��a��K<��|�k��^B��B�O@䮺>
p4/3���H§�S�ԴUa�SV�*ڇZ�s�=�Nea%BO��YQ�$��e��*��>� ��R0E�@-��=�E��up&�-�S}-7�Gм̀a���6- n���!�7�b4�3Bʫ���N�C��3��h&I<�HF�t������ ����I�[c�B��@A�
����t��qĬ��
{'71�C�^�f���Z��Ke�a�\�+`��ג���Z���Fw3��PIp� ��TY���G��g�˥)�o�zka6Ks>86�;38!���TX������0��e�����xI�e��<���43��S!.̀m�)$��i���#SOF̈́�ި�����F�51�[.���ȪIDQ}."���ESͿo��$rel�"� W��-�D>2f��X�DxD� \k�ϳ����t(�����P�
�Y3�0͙(j̆L*�� ���'����Y<�-!�ӑzx;3��?��s�-��g�������f������>����m�������=ݲ�M�(F�!�;3���	�u�j'�N�JE�1Of��oI,w;�0 �4΄}���VZ��x� ������s    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
.  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�͗mLSg�Ͻ���
���R�����!�s�eK\��dRP5ٟe&��f[����l�c�gqY�Mf��8�����!��R��BKKK���{�-���܏�����y�s�9��x���)��
 ðmH��B�|��V����n���]��hD�
<� 5�d0&xn��>��H��2��6;�$H��a�q��Z�D &[�N�/)*�]n�34�T&���d�����{��_�� >v٭�u}ssw5N���ڛ<48�8�F �ܖ �-�FL�[PX���7l�"d&X����.�� �)�,�¯��Ui4�L�v�2�����c̶���
��=�0�c>ڇ�Mߙ�kzYT�,5d���g�C��?�^?�)�����\A]��[�)T�9���{���%`�=)�Cjj:h�r� �@ܳN�Po0���n���w��i��I�y�3E� 'Jv�ե���s��]धX�c�����:��s��!� �6��rty���w&��v�@1r2! Z�O�Y���P�k��8x=�#,�-3��ч�5�+���mvՎ�RH)�y7�S������� ]r�B>_��Z��^��%���c�5sg�|�fg��;Hԅ��/����%�L��\D��[� �c�U���]�b�eY�y�*�E�����c�769��~�%��Ri8���m�Ji [�)�i�����^�����?�mu��{��HR���RM�Z�i�,�CW�h�U-	�������}ʔ����3~����^�!e�\�H�U0�g�dd�`+2z�
��#*o�	��+.ۯ%HRlO��
�P$�>k����SG�T�Z���#�+�U.fI)��� ���ٳ�	���+_��'o�j$��0�jZ	�����dI��ߌ���b�LF(	B�)� ����!�6m���������$���Ȗ�w�����0�d�A �x<�>$F���m�	�>��Ra�qM�@d-����oO
�8�B[�/9FKMR�Jl���XZ���f��� �m���2�?J�ޏ��j��Sc�}�D(�� ��� �!��0�督!	��{��Z`�9�22�U�2E�c|g���z�����[z^G��%M�?&���9��VW���ֶ@S��bcJZF�Ǳ����Hx
%���|������� �{J>�RrI�߮X�,1����FWQu�0�B���>� en�v5��
@���-I(����R�6�x>~f�P`8T5y�!f��$*8'�
@�؀
��e�!*)Pz}،����2�1���?��m��}�^�珂<���*v%���@\���oHG��E/��q���?º��kk�1XK�*�� 6
�K��~ �U�fR+@@�@�F֦9��p�����lH<y� ����h&٬    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�ŗoLgǿGK; �"L��S���W��:(m��2�E�\�Ө5ʌ�߂
�.ƨ�L&�&.���"�"Q0Q���B��F���m�{�ޕ�S�3I�������\�>w���0>dp����=dc��8 YN��Ҭ1�%�琳Y�Ť�gI	D1���HA�h��܎��vl��5�������\� ��%8RS���:���fU��Z477�#�o��	`Չ�--g� 
�0�n��	�� ͭα8
$� j�� ֜��Z[� �B�����-��S2@{�y6 �� �Du)�5��A��^��`�����ϧe��+�l �V��ªCjr|��r��e���"�9��߹Ý?o��{���Ł��G]3U K�C��H�=]��3bK٘#k�Pt�͚G�'�廓Sr�����	�{�
c��iaL@�ņAO��3��DR�����ᑵ�c�e4���� d��cpȯNl\9���Uw1��ϱ�) S7c�a4f�cj �d[1��4�N����!>ɘ�j����p8dc�0s�b̋-Z�̯���ͫ~2�S/���)��� ����4���	�˧geZ�׾�:��Fx�o_��9R�'b}�K,;��c�`4���1;�1# �hQö��?�2:����^ޏ�C�vmY"��՘NFc��SP ��*ґ ��S_iv�^��f@1�
����?vD��5�0�X����`4c�5n]��0�1�=]�� b�y�{3RS8�|��)]�R�� )�s`�o��K"��OP��s��`4c�u	*�0@�GF�1����t\�{�����1}� �V٘�
���yҧOJ2��YW�~O@fV�1���j;��F��5o����DZ<9Q��:�ă�kqD���Wٜ���ǖ�)TcVc��:y��DaM?W�a� DV�*�SL�'c&��������l̺����RN&9w����@pWM6R;֘o�3�ӵa����9�����ę��R�    IEND�B`�  Left(TopBitmap
         TPF0TEditorPreferencesDialogEditorPreferencesDialogLeft/Top� HelpType	htKeywordHelpKeywordui_editor_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionEditorPreferencesDialogClientHeight�ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxExternalEditorGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionC   Alternativ extern editor (påverkar bara redigering av fjärrfiler)TabOrder 	TCheckBoxExternalEditorTextCheckLeftTop-WidthQHeightCaptionH   Tvinga fram textöverföringsläge för filer redigerade i extern editorTabOrder  	TCheckBoxSDIExternalEditorCheckLeftTopWidthQHeightCaptionA   E&xtern editor öppnar varje fil i ett separat fönster (process)TabOrder    	TGroupBoxEditorGroup2LeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionEditorTabOrder 
DesignSize��   TRadioButtonEditorInternalButtonLeftTopWidth� HeightCaption&Intern editorTabOrder OnClickControlChange  TRadioButtonEditorExternalButtonLeftTop-Width� HeightCaption&Extern editorTabOrderOnClickControlChange  THistoryComboBoxExternalEditorEditLeft TopEWidthHeightAutoCompleteAnchorsakLeftakTopakRight TabOrderTextExternalEditorEditOnChangeControlChangeOnExitExternalEditorEditExit  TButtonExternalEditorBrowseButtonLeft1TopCWidthKHeightCaption   B&läddra...TabOrderOnClickExternalEditorBrowseButtonClick  TRadioButtonEditorOpenButtonLeftTopaWidth� HeightCaption&Associerad applikationTabOrderOnClickControlChange  TButtonDefaultButtonLeftTopxWidth� HeightCaption    Använd systemets standardeditorTabOrderOnClickDefaultButtonClick   	TGroupBox	MaskGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionAutomatiskt val av editorTabOrder
DesignSize�I  TLabel	MaskLabelLeftTopWidth� HeightCaption/   Använd den här editorn för &följande filer:FocusControlMaskEdit  THistoryComboBoxMaskEditLeftTop'WidthoHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder Text*.*OnExitMaskEditExit   TButtonOkButtonLeft� TopdWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� TopdWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft?TopdWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  	TCheckBoxRememberCheckLeftTopLWidthQHeightAnchorsakLeftakBottom Caption   &Kom ihåg den här editornTabOrder   TPF0TFileFindDialogFileFindDialogLeftoTop� HelpType	htKeywordHelpKeywordui_findBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionFindXClientHeight�ClientWidth2Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth�
ParentFont		Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                      '!�+$�PE;�th^���}������º�                                                                                                                                                                                                                                '!�+$�PE;�th^���}������º�����                                                                                                                                                                                                                            '!�+$�PE;�th^���}������º�����wg[�                                                                                                                                                                                                                        '!�+$�PE;�th^���}������º�����wg[�0("�                                                                                                                                                                                                                    '!�+$�PE;�th^���}������º�����wg[�0("�&!�                �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�        '!�+$�PE;�th^���}������º�����wg[�0("�&!�                    �vW����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������vW�    91)�.&!�PE;�th^���}������º�����wg[�0("�&!�                        �vW���������������������������������������������������������������������������������������������������������������������ô�������{n�yl`�yl`�{mb���u�����;���������������������������vW�ZK?�taS�m[N�tg]���}������º�����wg[�0("�&!�                            �vW�������������������������������������������������������������������������������������������������������������|oc�MA7�QD9�YK?�_PD�cRF�dTG�bRE�^OC�XI>�NA7�TH>��|p��ĵ�������������kWG�{i\��������xgY������º�����wg[�0("�&!�                                �vW�����������������������������������������������������������������������������������������������������dWL�OB8�`PD�n\N�r_Q�n[N�jXK�hWJ�gVI�hWJ�kYL�o\O�s`R�jYL�\MA�M@6�yl`��ȹ�����{i\������������������qd�����wg[�0("�&!�                                    �wX����������������������������������������������������������������������������������������������vj�NA7�bRE�r_Q�kZL�cRF�\MA�gYO��wn�������������sk�aSH�]NB�eTG�n\N�p^P�]NB�L@6�dTI�������������������������taS�2*$�&!�                                        �xY�����������������������������������������������������������������������������������������aUJ�VH=�o]O�lZM�_OC�vh]���������������������������������������������iZO�bRE�o]O�kYL�QD9�|rj���������������������taS�8/(�                                            �yY����������������������^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��vX�RD8�\MA�r_Q�dTG�iZO�������������������������������������������������������������`RF�iWJ�q^P�UG<�sjb�������������{i\�ZJ?�                                                �zZ���������������������������������������������������������������������������������_SH�]NB�q^P�`PD��uj���������������������������������������������������������������������qcW�eTG�r_Q�UG<�}sk�����{i\�[L@�                                                    �{Z�����������������������������������������������������������������������������|od�XJ>�r_Q�`PD���������������������������������������������������������������������������������xm�eTG�q^P�PC9�dUI�p^P�                                                        �{[�����������������������`���`���`���`���`���`���`���`���`���`���`���`���`��gO�PC8�q^P�cRF��uh��Ƿ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ��ʺ���������������������m^S�hWJ�kYL�J>4�I=1*                                                        �|\�������������������������������������������������������������������������WKA�gVI�jXK�m]R�����������������������������������������������������������������������������������������ɸ��_PD�o]O�]MB�K?4�                                                        �}\�������������������������������������������������������������������������TF;�r_Q�]NB�˽�������������������������������������������������������������������������������������������Ų�����bRE�p^P�M@6�G=46                                                    �~]�����������������������a���a���a���a���a���a���a���a���a���a���a���a�VG:�fUI�hWJ��sf��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű��ű����������������������ð�����eVK�n\N�\MA�K>5�                                                    �^������������������������������������������������������������������Ƚ�MA6�r_Q�_OC�Ŷ�����������������������������������������������������������������������������������������������¬���������dTG�kYL�K>5�@                                                  ��^���������������������������������������������������������������������XI>�o\O�\MB�������������������������������������������������������������������������������������������������������������]NB�s`R�OB7�K>5:                                                ��_�����������������������c���c���c���c���c���c���c���c���c���c���c�fSB�bRE�iXK��vg�������������������������������������������������������������������������������������������������׾����������bSH�o\O�WI=�J?4u                                                ��`�����������������������������������������������������������������bVL�hWJ�dTG�����������������������������������������������������������������������������������������������������׼����������{k_�kYL�^NC�J?5�                                                ��`�����������������������������������������������������������������VJ@�lZM�bRE�����������������������������������������������������������������������������������������������������׻�����������|m�iWJ�cRF�J>4�                                                ��a����������������������^��^��^��^��^��^��^��^��^��^��^�K?5�n\N�aQE�����Ը��ֽ��׿���������������������������������������������������������������������������������������������������p�gVI�eTH�J>5�                                                ��b�����������������������������������������������������������������RF<�lZM�aQE������������������������������������������������������������������������������������������������������«������׾��|l�hWJ�cSF�K?5�                                                ��b�����������������������������������������������������������������_TI�jXK�dSG������������������������������������������������������������������������������������������������������«������Թ�~l]�jYK�_PC�K?4�                                                ��c�����������������������`���`���`���`���`���`���`���`���`���`���`�aO?�dSG�hWJ��zh�Ե��׻���­��­��­��­��­��­��­��­��­��­��­��­��­��­��­��­��­����������������������Į������Թ�eUI�n\N�YJ?�K=3�                                                ��c���������������������������������������������������������������������ZK@�n[N�aRF��������������������������������������������������������������������������������������������������ű��ؿ��Ī�\MA�r_Q�PC9�H>4J                                                ��d�����������������������������������������������������������������ɾ��PC8�s`R�]NB�̸�����������������������������������������������������������������������������������������������Ű��պ�����bRF�n\N�K?5�@00                                                ��e�����������������������a���a���a���a���a���a���a���a���a���a���a���`�PC7�jYL�eUH��yh�ն��׻���ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ��ȵ���������������������پ���ҷ�m]P�kZL�`PD�J>4�                                                    ��f�������������������������������������������������������������������������XJ>�p^P�\MA�Ӿ������������������������������������������������������������������������������������������ظ������_OC�r_Q�OB8�H?2Q                                                    ��f�������������������������������������������������������������������������NB8�lZM�fUI�}k]�����������������������������������������������������������������������������������������ΰ��eTH�lZM�bRF�K>5�                                                       ��g�����������������������c���c���c���c���c���c���c���c���c���c���c���c���c�w_J�TF;�r_Q�_OC���o�ն��׹���ɷ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ��ͼ���������������������yfX�dTG�o]O�NA7�J<2L                                                        ��g�����������������������������������������������������������������������������dXN�`PD�o]O�]NB�����������������������������������������������������������������������������������s�`PD�r_Q�VH=�K?5�                                                            ��h���������������������������������������������������������������������������������RF<�fUH�n\N�]NB���s������������������������������������������������������������������ѽ��rb�`PD�q^P�\MA�K>5�I7$                                                            ��i�����������������������e���e���e���e���e���e���e���e���e���e���e���e���e���e���e��rW�M@5�fUH�o]O�_OC�~k\�¨��׷��׷��ټ���Į��˸��ξ������ξ��˹��Ű�ٽ��׷������ǳ��l[N�cRF�r_Q�]NB�K?5�K<5"                                                                ��i�������������������������������������������������������������������������������������ƾ��RF<�_PD�r_Q�fUI�\MA��|k�̸��������������������������������������į���rc�]NB�jYK�q^P�XI>�WH;�H;4'                                                                    ��j���������������������������������������������������������������������������������������������cXN�UG<�lZM�p]P�fUH�]NB�aRF��o����������������������wg�\MB�_OC�hWJ�r_Q�gVI�PC8�{pg���e�                                                                        ��k�����������������������g���g���g���g���g���g���g���g���g���g���g���g���g���g���g���g���g���g���e�yaL�L@5�XJ?�jYK�s`R�m[N�hWJ�dTG�bRE�bRE�bRE�eTH�iXK�o\O�r_Q�fUH�TF;�WLB�����������k�                                                                        ��k�������������������������������������������������������������������������������������������������������������UI?�PC8�[L@�cSF�iXK�lZM�n\O�lZM�hWJ�bRE�XJ>�MA6�`UL�������������������k�                                                                        ��l�������������������������������������������������������������������������������������������������������������������������xne�_TJ�PE;�K?5�UJ@�dYO�~sk�������������������������������l�                                                                        ��m�����������������������i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���i���k��Ϻ��κ��κ��κ��κ���m�                                                                        ��m������������������������������������������������������������������������������������������������������������������������������������������������������ǰ��ê��ê��ê��ê��ê��ê���m�                                                                        ��n����������������������������������������������������������������������������������������������������������������������������������������������ǰ�ҷ��ҷ��ҷ��ҷ��ҷ��ҷ��ҷ��ҷ����n�                                                                        ��o�����������������������k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���k���n���q���q���q���q���q�˫��˫��˫��˫��˫����o�                                                                        ��o���������������������������������������������������������������������������������������������������������������������������������ʪ��ßz�ßz�ßz�ßz�ßz�ßz�ßz�ßz�ßz�ßz�ßz���o�                                                                        ��p������������������������������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿���ª���p�                                                                        ��p�����������������������l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l��������������������������������������̹��ư�׿���ª���pԳ�f                                                                        ��q����������������������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿���ë���qԳ�f                                                                            ��r������������������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿���ë���rԿ�f                                                                                ��r�����������������������n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n��������������������������̹��ư�׿���ì���rԿ�f                                                                                    ��r����������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿���ì���rԿ�f                                                                                        ��r������������������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f                                                                                            ��r�����������������������p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p��������������̹��ư�׿��������rԿ�f                                                                                                ��r����������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f                                                                                                    ��r������������������������������������������������������������������������������������������������������������������������������̹��ư�׿��������rԿ�f                                                                                                        ��r������������������������������������������������������������������������������������������������������������������������������ư�׿��������rԿ�f                                                                                                            ��r�����������������������������������������������������������������������������������������������������������������������������׿��������rԿ�f                                                                                                                ��r�����������������������������������������������������������������������������������������������������������������������������������rҿ�f                                                                                                                    ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���rҿ�f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������� ������� ������� ������� �     0�      �      �      �      �      ?�      �      ��     ��     ��     ��     ��     ��     ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��     ��     ��     ��     ��     ��     ��     ��     ��     ?��     ?��     ?��     ?��     ?��     ?��     ?��     ?��     ?��     ?��     ?��     ��     ���    ���    ���    ���    ���    ���    ?���    ���    ����   ����   ���������������������������(   0   `          �%                                                                                                                                                                                              ' O-&�[PG��|s�����                                                                                                                                                                        ' O-&�[PG��|s�����Ƚ��                                                                                                                                                                    ' O-&�[PG��|s�����Ƚ���ym�                                                                                                                                                                ' O-&�[PG��|s�����Ƚ���ym�3+$�        �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�            ' O-&�[PG��|s�����Ƚ���ym�3+$�&!]        �vW����������������������������������������������������������������������������������������������������������������������������������vW�        ' O-&�[PG��|s�����Ƚ���ym�3+$�&!]            �vW����������������������������������������������������������������������������������������������������������������������������������vW�    ' O-&�[PG��|s�����Ƚ���ym�3+$�&!]                �vW����������������������������������������������������������������������������������������������Ǹ��ô������������������������������vW�PB8NB7�[PG��|s�����Ƚ���ym�3+$�&!]                    �wX����������������������������������������������������������������������������������th�SG<�K?5�K?5�K?5�K?5�MA7�uh]�����������������v^I��rf�����{j^�����Ƚ���ym�3+$�&!]                        �xY������������������^��^��^��^��^��^��^��^��^��^��^��^��~]�|bK�QC8�NB7�[MA�gVI�n\N�r_Q�s`R�o]O�iXK�^OC�RD:�MA7���z�Ƕ���sf���������������v��ym�3+$�&!]                            �yZ�����������������������������������������������������������������qdY�NA7�aQE�r_Q�vdX�����ĸ���ƽ�����Ƚ�������wj�r_Q�gVI�QD9�QD:���������������������QD:�&!]                                �zZ�������������������������������������������������������������_SH�TF;�o]O��nb�ʿ����������������������������������������}�q^P�ZL@�NB8��������������sg�L>5�                                    �{[�������������������`���`���`���`���`���`���`���`���`��{\�VG:�XJ>�q^P������ʼ���������������������������������������������ĸ��r_Q�`QD�NB8������rf�QD;�                                        �}\�����������������������������������������������������|od�SE:�q_Q��������������������������������������������������������������Ǽ�r_Q�[L@�PD9�hZHX                                            �~]�����������������������������������������������������L@6�n\N�������������������������������������������������������������������������q^P�QD9�J>4�                                            �^�������������������a���a���a���a���a���a���a���a�YJ<�\MA�saT�ҿ���Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ��Ǵ������������������ų���t�fUI�K?5�J55                                        ��_����������������������������������������������ʿ�K?5�o]O��������������������������������������������������������������������������ï�����r_Q�QD9�J?4q                                        ��`�������������������������������������������������TG<�p^P���������������������������������������������������������������������������������n`�^OC�J>5�                                        ��a�������������������c���c���c���c���c���c���c�aO?�`PD�wfY�������������������������������������������������������������������������ؿ����������jXK�K?5�@                                      ��a���������������������������������������������aUK�fUH��vh�������������������������������������������������������������������������׽������Ƴ��o\O�K?5�D<3                                    ��b���������������������������������������������PD:�iXK���r�������������������������������������������������������������������������ٿ������к��s`R�K?5�J;14                                    ��c�������������������e���e���e���e���e���e���e�QC8�hWJ��}m�غ���ì��ì��ì��ì��ì��ì��ì��ì��ì��ì��ì��ì��ì������������������«�����̴��r_Q�K?5�H=2.                                    ��d���������������������������������������������eYO�dTG��rb��������������������������������������������������������������������������í���������n\N�K?5�F:.                                    ��e���������������������������������������������{pf�]NB�q_Q��������������������������������������������������������������������������ư��׾���t�hWJ�K>5�                                        ��f�������������������g���g���g���g���g���g���g��jQ�QD9�r_Q�ĩ��ھ���ɴ��ɴ��ɴ��ɴ��ɴ��ɴ��ɴ��ɴ��ɴ��ɴ��ɴ��ɴ������������������Ű��ҷ�saR�[LA�J?4�                                        ��g�������������������������������������������������K?5�lZM���v���������������������������������������������������������������������ھ������r_Q�NB7�I>2[                                        ��h�������������������������������������������������zoe�WI>�p^P���������������������������������������������������������������������յ��zgX�bRE�J>5�333
                                        ��h�������������������i���i���i���i���i���i���i���i��~_�L?5�hWJ�~k[�Ҵ�������ν��Ͼ��Ͼ��Ͼ��Ͼ��Ͼ��Ͼ��Ͼ��Ͼ��Ͼ�������������������l�o]O�NA7�J>5o                                            ��i���������������������������������������������������������NA7�n\N��zj�������������������������������������������������������������q^P�SF;�K?5�@                                              ��j���������������������������������������������������������zof�RD:�n\N�|k[����������������������������������������������Ҿ���v�q_Q�WI>�K>4�I7.                                                ��k�������������������k���k���k���k���k���k���k���k���k���k���h�hUC�NA7�hWJ�p]P���u�Ū��ٹ��ں��۽��۾��ۻ��ں��̯������q`P�n\N�RE:�WH;�H;4'                                                    ��l���������������������������������������������������������������������L@6�WI>�lZM�r_Q�p^P��qa��}l���o��ue�weV�p^P�o]O�\MA�L@6�}rh���g�                                                        ��m�������������������������������������������������������������������������|rj�K?5�QD9�]NB�dSG�hWJ�iWJ�eTH�_PD�TG<�K?5�f[P�����������m�                                                        ��n�������������������l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���e��oU�kWE�\L=�QD8�OB7�YJ<�eSB��iQ�¯���ɳ��ɳ��ɳ���n�                                                        ��o���������������������������������������������������������������������������������������������������������׾��Ҷ��Ҷ��Ҷ��Ҷ��Ҷ����o�                                                        ��o�������������������������������������������������������������������������������������������������ҷ��ţ�ţ�ţ�ţ�ţ�ţ�ţ���o�                                                        ��p�������������������n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n���n������������������������������Ͻ��Ȳ�ּ����p�                                                        ��q������������������������������������������������������������������������������������������������������������������Ͻ��Ȳ�ֽ����q���U                                                        ��r��������������������������������������������������������������������������������������������������������������Ͻ��Ǳ�־����q���U                                                            ��r�������������������p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p������������������Ͻ��Ǳ�־����q���U                                                                ��r������������������������������������������������������������������������������������������������������Ͻ��Ǳ�־����q���U                                                                    ��r��������������������������������������������������������������������������������������������������Ͻ��Ǳ�־����q���U                                                                        ��r����������������������������������������������������������������������������������������������Ͻ��Ǳ�׾����q���U                                                                            ��r����������������������������������������������������������������������������������������������Ǳ�׾����q���U                                                                                ��r���������������������������������������������������������������������������������������������׾����q���U                                                                                    ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���q���U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������  ������  ������  �����   �      �     �     �      �      �      �    ?  �      �    �  �   �  �   �  �    �  �    �  �    �  �      �      �      �      �      �    �  �    �  �    �  �    �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   ?�  �   �  �   ��  �  ��  �  ��  �  ��  �  ��  ������  ������  (   (   P          @                                                                                                                                                          #:' �>4,�dVL�}od���{�                                                                                                                                    #:' �>4,�dVL�}od���{���x�                                                                                                                                #:' �>4,�dVL�}od���{���x�,& �    �wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX��wX�#:' �>4,�dVL�}od���{���x�,& �&!]    �xY������������������������������������������������������������������������������������������������������������������dK�' �>4,�dVL�}od���{���x�,& �&!]        �yZ������������������������������������������������������������������������������Ƹ�;������������������������������8/'�>4,�dVL�}od���{���x�,& �&!]            �zZ��������������������������������������������������������������Ⱥ���v�]QF�OB8�VH=�YK?�RE:�OC9�xl`����������´�q_Q�����}qg�}od���{���x�,& �&!]                �{[����������������������������������������������������������xl�PC9�p^Q��sc���o���z������r��|j�|hY�\MA�]QF�kZM�������������������x�,& �&!]                    �}\��������������������������������������������������ɼ�^RG�jYL��|k�ò���������������������������ƻ���~��l\�QD9�������������Ż��8/(�&!]                        �~]���������������p���p���p���p���p���p���p���p���h�QD8�zgX������˻�������������������������������������Ǵ���yh�XJ?������ž�wdW�SF<�                            �^���������������������������������������������eXN�ubT������������������������������������������������������ʾ��zi�RE:�hWK�bQFu                                ��_���������������������������������������������aQE�������������������������������������������������������������ͼ���o_�M@6�@                                  ��`���������������p���p���p���p���p���p���l�PC7��wf�ҽ���ι��ι��ι��ι��ι��ι��ι��ι��ι��ι��ι��ι��ι�������������_PD�I?4v                                ��a�����������������������������������������^OC����������������������������������������������������������������������Ĵ��n^�K?5�                                ��a��������������������������������������zp�vdU�͹�����������������������������������������������������������������������~m�MA7�J55                            ��b���������������p���p���p���p���p���p�aP@��qa�Ӻ���Ū��Ū��Ū��Ƭ��ǭ��Ȯ��ȯ��ȯ��ȯ��ȯ��ȯ��Ǯ��Ƭ��ƫ���������������z�XJ?�H<3<                            ��c�������������������������������������]QG��wf��н�������������������������������������������������������������������������`PD�K>5R                            ��d�������������������������������������_TJ��ud��͹�����������������������������������������������������������������������~�^OC�I=3P                            ��e���������������p���p���p���p���p���p�cQA��n^�д���ũ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ��ʲ���������������u�VI=�G=46                            ��f���������������������������������������~�p^P�Ĭ�������������������������������������������������������������������Ѽ��{j�J>4�@++                            ��g�����������������������������������������XJ?���y�����������������������������������������������������������������ζ��|hY�J>5�                                ��h���������������p���p���p���p���p���p���o�YJ<��n^�ɭ�������м��н��н��н��н��н��н��н��н��н��н��н�����������s�WI>�I=4T                                ��h���������������������������������������������XJ>���p��͸���������������������������������������������������������wdV�K?5�                                   ��i����������������������������������������������vl�fUI���z��Ϻ���������������������������������������������ī���qa�QC8�I>41                                    ��j���������������p���p���p���p���p���p���p���p���m�^N?�gVI���p�˯��ݾ���ƫ��θ��Ҿ������м��˳�����ո�������n^�PC9��tX�                                        ��k�����������������������������������������������������~sj�ZL@��p`���}�̴���ʵ����������ϻ�ֿ�������|k�n]O�VJ@��û���k�                                        ��l�������������������������������������������������������������\QG�\NB�vcU��sc��{i��}l��wf��l\�iXK�OC8��|s�����������l�                                        ��m���������������p���p���p���p���p���p���p���p���p���p���p���p���n��x[�r]I�ZJ<�NB7�K?5�TF:�fTC��kS���g���������������m�                                        ��n����������������������������������������������������������������������������������������������ʴ��ɲ��ɲ��ɲ��ɲ���n�                                        ��o�����������������������������������������������������������������������������������������Ҷ��Ҷ��Ҷ��Ҷ��Ҷ��Ҷ����o�                                        ��o���������������p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p������������������������������ɴ�Լ����o�                                        ��p������������������������������������������������������������������������������������������������������ɴ�ּ����p���U                                        ��q��������������������������������������������������������������������������������������������������ȳ�ֽ����q���U                                            ��r���������������p���p���p���p���p���p���p���p���p���p���p���p���p���p���p���p������������������ȳ�־����q���U                                                ��r������������������������������������������������������������������������������������������ȳ�־����q���U                                                    ��r��������������������������������������������������������������������������������������ȳ�־����q���U                                                        ��r����������������������������������������������������������������������������������ȳ�־����q���U                                                            ��r���������������������������������������������������������������������������������׾����q���U                                                                ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���q���U                                                                                                                                                                                                                                �����   �����   ����    �       �      �      �      �      �      �   ?   �      �      �      �      �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �      �      �      �   �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  ?�   �  �   �  ��   �����   (       @          �                                                                                                                                      &!�4,%�`SH�                                                                                                                &!�4,%�`SH��rf�                                                                                                            &!�4,%�`SH��rf�����    �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�        &!�4,%�`SH��rf�����[QI�    �vW������������������������������������������������������������������ĵ��ô��������������vW�   F;2�4,%�`SH��rf�����[QI�&!�    �wX���������������������������������������������������������eXM�\MA�eUH�fUI�^OC�_SH���z��qT�cTGÛ��������rf�����[QI�&!�        �xY�������������������������������������������������YLA�vcU���|�ѿ�����������µ�����{gX�UG<�tg\�������������[QI�&!�            �zZ��������������yY��yY��yY��yY��yY��yY��yY�x^H�]NB���y�κ���´��õ��õ��õ��õ�������������dTH���}���������B8/�                �|[�������������������������������������µ��[MA�������������������������������������������������cSG�vg]�aPE�                    �}]��������������|\��|\��|\��|\��|\��z[�VH:���s�Ѽ��ӿ��ӿ��ӿ��ӿ��ӿ��ӿ��ӿ��������������Ӿ������SF:�J55                    �^�������������������������������������q_Q�������������������������������������������������ӽ������zgX�J>5�                    ��_��������������^��^��^��^��^�`N>��}l�ҹ��ҹ��ҹ��ҹ��ҹ��ҹ��ҹ��ҹ��ҹ��������������Ӻ��������x�M@6�                    ��a���������������������������������UG<�«��������������������������������������������������ҷ������¬��\MA�I7.                ��b���������������a���a���a���a��~]�[LA�Ȯ��ӷ�������ư��˷��˷��˷��˷��˷��˷���������������������ͷ��dTG�J;14                ��c���������������������������������ZL@�θ���������������������������������������������������ѿ�����˲��cTG�G=32                ��e���������������c���c���c���c���c�SE:�����׻����������������������������������������������������������ZL@�@33                ��f���������������������������������{pf��ud�����������������������������������������������������������p�J?4�                    ��g���������������f���f���f���f���f��mS�jZL�ϲ���ǯ���������������������������������������������պ��taS�J>4                    ��h�������������������������������������h[R��zi���������������������������������������������ֶ����o�PC9�I7$                    ��j���������������h���h���h���h���h���h��}^�XJ>���x�Է���̷�����������������������������������y�[L@�J=4S                        ��k�����������������������������������������ú��YK@��zi��Ʊ��������������������������̷���r�ZK@�K=4p                            ��l���������������k���k���k���k���k���k���k���k��`�]M?�jYL��sc�����̱��β��¨���xg�o]P�WI;�I?5M                                ��n���������������������������������������������������������um�VI?�ZK@�ZL@�TG;�o`Q���u���l�                                    ��o���������������m���m���m���m���m���m���m���m���m���m���m���������ĥ����}�ǥ��ǥ��ǥ����o�                                    ��p������������������������������������������������������������������������������̸��ª���p�                                    ��q���������������p���p���p���p���p���p���p���p���p���p���p������������������̸��«���qҳ�f                                    ��r����������������������������������������������������������������������̸��ë���rɿ�f                                        ��r������������������������������������������������������������������̸��ë���rſ�j                                            ��r��������������������������������������������������������������̸�������rſ�j                                                ��r�������������������������������������������������������������������rſ�j                                                    ��r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���r���rÿ�j                                                                                                                                                                                    �������������  ��   �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?�  �  ��  ��  ��  �� �� �� �� �� �����(      0          `	                                                                                                     & �@7/��rf�    �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�   & �@7/��rf�}pf�    �vW��������������������������������������������������ȹ��������������sU�;2+�@7/��rf�}pf�'"�    �wX�����������������������������������������eXM�`QD�gWJ�bSF�^QE�����p\L�����}qg�}pf�'"�       �yZ����������^��^��^��^��^��|\�bP@�o]P�����ı��ʸ��ƴ������yfW�UH<���������<2+�           �{[�����������������������������~qf�|hY�Ͽ���������������������������yh�TG<�fUI�..            �~]�����������a���a���a���a��nS�iXK�­���ɷ��ɷ��ɷ��ɷ��ɷ���������ͺ��yfW�J?3�                ��_�������������������������}qg��yh����������������������������������î�����OB8�               ��`�����������c���c���c���c�XI=�����ٿ��ٿ��������������������������ؾ��̸��aQE�H80             ��b�������������������������ZL@�������������������������������������ؾ��Ի��fVI�H=2.            ��d�����������f���f���f���f�YJ<���|�ڽ���Ű��Ű��Ű��Ű��Ű���������ٿ��Ī��_PD�E;1            ��e���������������������������v��qa���������������������������������ټ����t�MA5�                ��g�����������h���h���h���h��}^�]NB�����۾���ν��Ͼ��Ͼ��Ͼ�������������n\O�J>4g                ��i���������������������������������kZM�������������������������Ŭ��{gX�K>5�                   ��j�����������k���k���k���k���k���j�}eN�^OC��p`���}����������xg�gWJ�mXF�@++                    ��l�������������������������������������������{�cWN�YK@�_QG�zk]�������l�                        ��n�����������m���m���m���m���m���m���m���m���������г��ɩ��ɩ��ɩ����n�                        ��p����������������������������������������������������������ϼ�������p�                        ��q�����������p���p���p���p���p���p���p���p��������������ϼ��«���qҳ�f                        ��r��������������������������������������������������ϼ��ë���rſ�j                            ��r����������������������������������������������ϼ��ª���rſ�j                                ��r���������������������������������������������׿����rſ�j                                    ��r���r���r���r���r���r���r���r���r���r���r���r���rÿ�j                                                                                                                                    ��� �   �   �   �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � ? �  � � �� ��� (      (          �                                                                                      $!M4,$�yk`��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�    $!M4,$�yk`�sg^��wX������������������������������������������������������wX�5/'\4,$�yk`�sg^�' v�xY�������������������������������������ocX�]QF�ocX������jR��wi�uh^�sg^�' v    �zZ�������w���w���w���w���w���h�VH<���������������������PC8���������9/(�        �|[�������������������������ZND��������������������������µ�L@6�bRF�            �}]�������w���w���w���w�zdR������ɶ��ɶ��ɶ��ɶ��ɶ�����Կ������J>5�            �^���������������������bVM�����������������������������Ӻ������K>5�            ��_�������}���}���}���}�L?5��©��˶��о������������������¬�����K?5�            ��a���������������������]QG����������������������������������ж�K>4�            ��b���������������������vcQ�γ������������������������������ë��J>4�            ��c�������������������������h[O�������������������������ֹ��VI>�J</&            ��d�����ť��ť��ť��ť��ť����l�jYL�Ӹ���ʲ��ѽ��ʲ��î�\NB�I>5W                ��f����������������������������������zr�QF<�l]Q�PC9�saO��{]�                    ��g�����ʪ��ʪ��ʪ��ʪ��ʪ��ʪ��ʪ����������������r���r���g�                    ��h��������������������������������������������������ʸ���g�                    ��j����������������������������������������������ʸ���j˳�f                    ��k������������������������������������������ɶ���jŪ�j                        ��l���l���l���l���l���l���l���l���l���l���l���kŪ�j                                                                                                            ���             0   p   p   p   p   p   p   p   �  �  �  �  �  �  � ��� (                 @                  �vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW��vW�    #:4+$�pe��xX������������������������������������������xX�#:4+$�pe�\QI��{[���������������������ö��ui^�TG=�TG=�ui^��iO�m_T�}nc�\QI�#:�~]�������h���h���h�|dM�vkb�����������������vja��|s��~u�#:    ��`�������������ø��ymd�������������������������pf]�RD:        ��b�������h���h�dRA������������������������������ǻ�K?4�        ��d�������������SG=��������������������������Ҽ�����K?4�        ��g�������k���k�PC7��˰�����������������������������K?4�        ��i�������������wlc��İ�������������������������и��J>5�        ��l�������m���m��z\�raR��ʹ������������������Ϸ�n_P�I?4I        ��n���������������������wi[��Ű���������Ӻ��scS�J>5�            ��q�������p���p���p���p��|_�{ri�TH>�SG<�qbT��y]�                ��r����������������������������������«���rͿ�f                ��r������������������������������ª���rſ�j                    ��r���r���r���r���r���r���r���r���rſ�j                                                                                                                                     ?  ��  
KeyPreview	OldCreateOrderPositionpoOwnerFormCenterOnClose	FormCloseOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize2� PixelsPerInch`
TextHeight 	TGroupBoxFilterGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionFilterTabOrder 
DesignSize�  TLabel	MaskLabelLeft1TopWidth/HeightCaption	&Filmask:FocusControlMaskEdit  TLabelRemoteDirectoryLabelLeft1TopGWidth0HeightCaption   Sö&k i:FocusControlRemoteDirectoryEdit  	TPaintBoxAnimationPaintBoxLeftTopWidth Height   THistoryComboBoxRemoteDirectoryEditLeft1TopWWidthvHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxMaskEditLeft1Top$Width HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextMaskEditOnChangeControlChangeOnExitMaskEditExit  TStaticTextMaskHintTextLeft� Top;Width|Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	  TButton
MaskButtonLeftWTop"WidthPHeightAnchorsakTopakRight Caption	&RedigeraTabOrderOnClickMaskButtonClick   TButtonStartStopButtonLeft�TopWidthlHeightAnchorsakTopakRight Caption&StartXDefault	TabOrderOnClickStartStopButtonClick  TButton
HelpButtonLeft�Top*WidthlHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TIEListViewFileViewLeftTop� Width�Height� AnchorsakLeftakTopakRightakBottom FullDrag	ReadOnly		RowSelect		PopupMenuFileViewPopupMenuTabOrder	ViewStylevsReport
OnDblClickFileViewDblClickOnEnterControlChangeOnExitControlChange
NortonLikenlOffColumnsCaptionNamnWidthP CaptionKatalogWidthx 	AlignmenttaRightJustifyCaptionStorlekWidthP Caption   ÄndradWidthZ  	OnCompareFileViewCompareOnContextPopupFileViewContextPopupOnSelectItemFileViewSelectItem  
TStatusBar	StatusBarLeft Top�Width2HeightPanels SimplePanel	  TButtonFocusButtonLeft�Top� WidthlHeightActionFocusActionAnchorsakTopakRight TabOrder  TButton
CopyButtonLeft�TopqWidthjHeightAction
CopyActionAnchorsakRightakBottom TabOrder  TButtonDeleteButtonLeft�Top� WidthlHeightActionDeleteActionAnchorsakTopakRight TabOrder  TButtonDownloadButtonLeft�Top� WidthlHeightActionDownloadActionAnchorsakTopakRight TabOrder  TButton
EditButtonLeft�Top� WidthlHeightAction
EditActionAnchorsakTopakRight Caption	&RedigeraTabOrder  
TPopupMenuFileViewPopupMenuLeft�Top 	TMenuItemFocus1ActionFocusActionDefault	  	TMenuItemN1Caption-  	TMenuItemEdit1Action
EditAction  	TMenuItem	Download1ActionDownloadAction  	TMenuItemDelete1ActionDeleteAction  	TMenuItemN2Caption-  	TMenuItemSelectAllItemActionSelectAllAction  	TMenuItemN3Caption-  	TMenuItemCopyResults1Action
CopyAction   TActionList
ActionListLeft�Top= TActionDeleteActionCaption&Ta bortSecondaryShortCuts.StringsF8 ShortCut.	OnExecuteDeleteActionExecute  TActionFocusActionCaptionF&okus	OnExecuteFocusActionExecute  TActionSelectAllActionCaptionM&arkera alltShortCutA@	OnExecuteSelectAllActionExecute  TAction
CopyActionCaption&Kopiera resultatShortCutC@	OnExecuteCopyActionExecute  TActionDownloadActionCaptionLadda &ner...ShortCutt	OnExecuteDownloadActionExecute  TAction
EditActionCaption	&RedigeraSecondaryShortCuts.StringsCtrl+E ShortCuts	OnExecuteEditActionExecute      TPF0TFileSystemInfoDialogFileSystemInfoDialogLeft@Top� HelpType	htKeywordHelpKeyword	ui_fsinfoBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption#Information om server och protokollClientHeight�ClientWidthsColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSizes� PixelsPerInch`
TextHeight TButtonCloseButtonLeft� ToplWidthKHeightAnchorsakRightakBottom Cancel	Caption   StängDefault	ModalResultTabOrder  TButton
HelpButtonLeftToplWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPageControlPageControlLeft Top WidthsHeight`
ActivePageProtocolSheetAlignalTopAnchorsakLeftakTopakRightakBottom TabOrder OnChangePageControlChange 	TTabSheetProtocolSheetCaption	Protokoll
DesignSizekD  	TGroupBoxHostKeyGroupLeftTop� Width_HeightWAnchorsakLeftakRightakBottom Caption$   Nyckelfingeravtryck till värdserverTabOrder
DesignSize_W  TLabelLabel2Left
TopWidth1HeightCaptionAlgoritmFocusControlHostKeyAlgorithmEdit  TLabelLabel3Left
Top)Width.HeightCaptionSHA-256:FocusControlHostKeyFingerprintSHA256Edit  TLabelLabel4Left
Top@WidthHeightCaptionMD5:FocusControlHostKeyFingerprintMD5Edit  TEditHostKeyFingerprintSHA256EditLeftATop)WidthHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFace	PopupMenuFingerprintPopupMenuReadOnly	TabOrderTextHostKeyFingerprintSHA256EditOnContextPopup(HostKeyFingerprintSHA256EditContextPopup  TEditHostKeyAlgorithmEditLeftATopWidthHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextHostKeyAlgorithmEdit  TEditHostKeyFingerprintMD5EditLeftATop@WidthHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFace	PopupMenuFingerprintPopupMenuReadOnly	TabOrderTextHostKeyFingerprintMD5EditOnContextPopup(HostKeyFingerprintSHA256EditContextPopup   	TListView
ServerViewLeftTopWidth_Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�  Caption   VärdeWidth�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup  	TGroupBoxCertificateGroupLeftTop&Width_HeighthAnchorsakLeftakRightakBottom CaptionCertifikatets fingeravtryckTabOrder
DesignSize_h  TLabelLabel5Left
TopWidth.HeightCaptionSHA-256:FocusControl CertificateFingerprintSha256Edit  TLabelLabel6Left
Top+Width"HeightCaptionSHA-1:FocusControlCertificateFingerprintSha1Edit  TEdit CertificateFingerprintSha256EditLeftATopWidthHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder Text CertificateFingerprintSha256Edit  TButtonCertificateViewButtonLeft
TopBWidthyHeightCaption   &Fullständigt certifikatTabOrderOnClickCertificateViewButtonClick  TEditCertificateFingerprintSha1EditLeftATop+WidthHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFace	PopupMenuFingerprintPopupMenuReadOnly	TabOrderTextCertificateFingerprintSha1EditOnContextPopup(HostKeyFingerprintSHA256EditContextPopup    	TTabSheetCapabilitiesSheetCaption   Möjligheter
ImageIndex
DesignSizekD  	TGroupBox	InfoGroupLeftTop� Width_HeightrAnchorsakLeftakRightakBottom Caption   Övrig informationTabOrder
DesignSize_r  TMemoInfoMemoLeft	TopWidthMHeightWTabStopAnchorsakLeftakTopakRight 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneColor	clBtnFaceLines.StringsInfoMemo 
ScrollBarsssBothTabOrder WordWrap   	TListViewProtocolViewLeftTopWidth_Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�  Caption   VärdeWidth�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup   	TTabSheetSpaceAvailableSheetCaption   Tillgängligt utrymme
ImageIndex
DesignSizekD  TLabelLabel1LeftTopWidthHeightCaption
   &Sökväg:FocusControlSpaceAvailablePathEdit  	TListViewSpaceAvailableViewLeftTop(Width_Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�  Caption   VärdeWidth�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupControlContextPopupOnCustomDrawItem SpaceAvailableViewCustomDrawItem  TEditSpaceAvailablePathEditLeft8Top	Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnEnterSpaceAvailablePathEditEnterOnExitSpaceAvailablePathEditExit  TButtonSpaceAvailableButtonLeft TopWidthcHeightAnchorsakTopakRight CaptionKon&trolleraTabOrderOnClickSpaceAvailableButtonClick    TButtonClipboardButtonLeftToplWidth� HeightAnchorsakRightakBottom Caption&Kopiera till urklippTabOrderOnClickClipboardButtonClick  
TPopupMenuListViewMenuLeft� Topb 	TMenuItemCopyCaptionK&opieraOnClick	CopyClick   
TPopupMenuFingerprintPopupMenuLeft� Topb 	TMenuItemCopy1ActionEditCopyAction  	TMenuItem ActionEditSelectAllAction   TActionListFingerprintActionListLeftHTopb 	TEditCopyEditCopyActionCategoryEditCaptionK&opieraShortCutC@	OnExecuteEditCopyActionExecuteOnUpdateEditCopyActionUpdate  TEditSelectAllEditSelectAllActionCategoryEditCaption&Markera alltShortCutA@     TPF0TFullSynchronizeDialogFullSynchronizeDialogLeftmTop� HelpType	htKeywordHelpKeywordui_synchronizeBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynkroniseraClientHeight�ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize�w  TLabelLocalDirectoryLabelLeft1TopWidthJHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft1TopDWidthWHeightCaption   F&järrka&talog:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  THistoryComboBoxRemoteDirectoryEditLeft1TopTWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeft1Top#WidthBHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeftzTop!WidthKHeightAnchorsakTopakRight Caption   Bl&äddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButtonOkButtonLeft� Top�WidthXHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrderOnClickOkButtonClickOnDropDownClickOkButtonDropDownClick  TButtonCancelButtonLeft;Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder	  	TGroupBoxOptionsGroupLeftTop� Width/HeightaCaption   Alternativ för synkroniseringTabOrder
DesignSize/a  	TCheckBoxSynchronizeDeleteCheckLeftTopWidth� HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top,Width� HeightAnchorsakLeftakTopakRight CaptionBara &valda filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight Caption&Endast existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizePreviewChangesCheckLeftTop,Width� HeightCaption   Fö&rhandsvisa ändringarTabOrderOnClickControlChange   TButtonTransferSettingsButtonLeftTop�Width� HeightAnchorsakLeftakBottom Caption   Överf&öringsinställningar...TabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxDirectionGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight Caption   Riktning/målkatalogTabOrder TRadioButtonSynchronizeBothButtonLeftTopWidth� HeightCaption   &BådaChecked	TabOrder OnClickControlChange  TRadioButtonSynchronizeRemoteButtonLeft� TopWidth� HeightCaption   &FjärrTabOrderOnClickControlChange  TRadioButtonSynchronizeLocalButtonLeft0TopWidth� HeightCaption&LokalTabOrderOnClickControlChange   	TGroupBoxCompareCriterionsGroupLeft=Top� Width� HeightaAnchorsakLeftakTopakRight Caption   JämförelsekriterierTabOrder
DesignSize� a  	TCheckBoxSynchronizeByTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Ä&ndringstidTabOrder OnClickControlChange  	TCheckBoxSynchronizeBySizeCheckLeftTop,Width� HeightAnchorsakLeftakTopakRight CaptionF&ilstorlekTabOrderOnClickControlChange  	TCheckBoxSynchronizeCaseSensitiveCheckLeftTopDWidth� HeightAnchorsakLeftakTopakRight Caption   Sk&riftlägeskänsligTabOrderOnClickControlChange   	TCheckBoxSaveSettingsCheckLeftTopUWidth�HeightAnchorsakLeftakTopakRight Caption   Använd &samma val nästa gångTabOrder  	TGroupBoxCopyParamGroupLeftTopjWidth�Height2AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamGroupClick   TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrder
OnClickHelpButtonClick  	TGroupBox	ModeGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight CaptionMetodTabOrder TRadioButtonSynchronizeFilesButtonLeftTopWidth� HeightCaptionSynkronisera &filerTabOrder OnClickControlChange  TRadioButtonMirrorFilesButtonLeft� TopWidth� HeightCaptionS&pegelfilerTabOrderOnClickControlChange  TRadioButtonSynchronizeTimestampsButtonLeft0TopWidth� HeightCaption   Synkronisera tidss&tämplarTabOrderOnClickControlChange   
TPopupMenuOkMenuLeft�Toph 	TMenuItemStart1Caption&StartDefault	OnClickStart1Click  	TMenuItemStartInNewWindowItemCaption   Starta i &nytt fönsterOnClickStartInNewWindowItemClick    TPF0TGenerateUrlDialogGenerateUrlDialogLeftqTopHelpType	htKeywordHelpKeywordui_generateurlBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionGenerate URL XClientHeightRClientWidth�Color	clBtnFaceConstraints.MinHeight,Constraints.MinWidth�
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize�R PixelsPerInch`
TextHeight TPageControlOptionsPageControlLeftTopWidth�Heighto
ActivePageUrlSheetAnchorsakLeftakTopakRight TabOrder OnChangeControlChange 	TTabSheetUrlSheetCaptionURL 	TCheckBoxUserNameCheckTagLeftTopWidth� HeightCaption   &AnvändarnamnTabOrder OnClickControlChange  	TCheckBoxHostKeyCheckTagLeft� TopWidth� HeightCaption   SSH &värdnyckelTabOrderOnClickControlChange  	TCheckBoxWinSCPSpecificCheckTagLeft� TopWidth� HeightCaptionWinSCP-specifikTabOrderOnClickControlChange  	TCheckBoxSaveExtensionCheckTag Left� Top6Width� HeightCaption   &Spara sessionsinställningarTabOrderOnClickControlChange  	TCheckBoxRemoteDirectoryCheckTagLeftTop6Width� HeightCaptionInitial &katalogTabOrderOnClickControlChange  	TCheckBoxPasswordCheckTagLeftTopWidth� HeightHelpType	htKeywordCaption
   &LösenordTabOrderOnClickControlChange  	TCheckBoxRawSettingsCheckTag@Left7TopWidth� HeightCaption   &Avancerade inställningarTabOrderOnClickControlChange   	TTabSheetScriptSheetCaptionSkript
ImageIndex TLabelLabel2LeftTopWidth&HeightCaption&Format:FocusControlScriptFormatCombo  TLabelScriptDescriptionLabelLeftTop Width�Height*AutoSizeCaptionScriptDescriptionLabelShowAccelCharWordWrap	  	TComboBoxScriptFormatComboLeftpTopWidthyHeightStylecsDropDownListTabOrder OnChangeControlChangeItems.Strings	SkriptfilBatchfilKommandoradPowerShell-skript    	TTabSheetAssemblySheetCaption.NET assemblerkod
ImageIndex TLabelLabel1LeftTopWidth3HeightCaption   &SpråkFocusControlAssemblyLanguageCombo  TLabelAssemblyDescriptionLabelLeftTop Width�Height*AutoSizeCaptionAssemblyDescriptionLabelShowAccelCharWordWrap	  	TComboBoxAssemblyLanguageComboLeftpTopWidthyHeightStylecsDropDownListTabOrder OnChangeControlChangeItems.StringsC#VB.NET
PowerShell     	TGroupBoxResultGroupLeftTopzWidth�Height� AnchorsakLeftakTopakRightakBottom CaptionResultXTabOrder
DesignSize��   TMemo
ResultMemoLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneTabOrder    TButton	CancelBtnLeft>Top1WidthKHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  TButton
HelpButtonLeft�Top1WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClipboardButtonLeftTop1Width� HeightAnchorsakLeftakBottom Caption&Kopiera till urklippTabOrderOnClickClipboardButtonClick   TPF0TImportSessionsDialogImportSessionsDialogLeftjTop� HelpType	htKeywordHelpKeyword	ui_importBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionImport sitesXClientHeightClientWidthwColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSizew PixelsPerInch`
TextHeight TLabelLabelLeftTopWidth=HeightCaption   &Importera från:FocusControlSourceComboBox  TButtonOKButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  	TListViewSessionListView2LeftTop'WidthiHeight� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsWidth�   ColumnClickDoubleBuffered	HideSelectionReadOnly	ParentDoubleBufferedParentShowHintShowColumnHeadersShowHint	TabOrder	ViewStylevsReport	OnInfoTipSessionListView2InfoTipOnKeyUpSessionListView2KeyUpOnMouseDownSessionListView2MouseDown  TButtonCheckAllButtonLeftTop� WidthqHeightAnchorsakLeftakBottom CaptionMarkera/avmarkera &allaTabOrderOnClickCheckAllButtonClick  TButton
HelpButtonLeft&Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  	TComboBoxSourceComboBoxLeftjTop
WidthxHeightStylecsDropDownListTabOrder OnSelectSourceComboBoxSelectItems.StringsPuTTY	FileZillaknown_hosts   TPanel
ErrorPanelLeft0Top\WidthHeighta
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder TLabel
ErrorLabelLeft Top WidthHeightaAlignalClient	AlignmenttaCenterCaption
ErrorLabelShowAccelCharLayouttlCenterWordWrap	   TButtonPasteButtonLeft� TopWidthKHeightCaptionKl&istra inTabOrderOnClickPasteButtonClick      TPF0TLicenseDialogLicenseDialogLeft�Top� ActiveControlCloseButtonBorderIconsbiSystemMenu BorderStylebsDialogCaption   AnvändarlicensClientHeight@ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenter
DesignSize�@ PixelsPerInch`
TextHeight TButtonCloseButtonLeft�TopWidthKHeightAnchorsakRightakBottom Cancel	Caption   StängDefault	ModalResultTabOrder   TMemoLicenseMemoLeftTopWidth�HeightAnchorsakLeftakTopakRight Color	clBtnFaceReadOnly	
ScrollBars
ssVerticalTabOrderWantReturns      TPF0TLocationProfilesDialogLocationProfilesDialogLeftWTop� HelpType	htKeywordHelpKeywordui_locationprofileBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionPlatsprofilerClientHeight�ClientWidth-Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize-� PixelsPerInch`
TextHeight TLabelLocalDirectoryLabelLeft.TopWidthJHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft.Top8WidthWHeightCaption   F&järrkatalog:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  TButtonOKBtnLeft/Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTophWidthHeight 
ActivePageSessionProfilesSheetAnchorsakLeftakTopakRightakBottom TabOrder 	TTabSheetSessionProfilesSheetTagCaptionSessionsplatsprofiler
DesignSize  	TTreeViewSessionProfilesViewTagLeft
Top	Width�Height� AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentParentDoubleBufferedTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDragItems.NodeData
                ��������           1 "           ��������            1 1             ��������            2             ��������            3            ��������           4 "           ��������            4 1             ��������            5   TButtonAddSessionBookmarkButtonTagLeft�Top	WidthSHeightAnchorsakTopakRight Caption   &Lägg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeft�Top)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�Left�Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonRenameSessionBookmarkButtonTagLeft�TopIWidthSHeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSessionBookmarkMoveToButtonTagLeft�TopiWidthSHeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick   	TTabSheetSharedProfilesSheetTagCaptionDelade platsprofiler
ImageIndex
DesignSize  	TTreeViewSharedProfilesViewTagLeft
Top	Width�Height� AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentParentDoubleBufferedTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDragItems.NodeData
                ��������           1 "           ��������            1 1             ��������            2             ��������            3            ��������           4 "           ��������            4 1             ��������            5   TButtonAddSharedBookmarkButtonTagLeft�Top	WidthSHeightAnchorsakTopakRight Caption   &Lägg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeft�Top)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonRenameSharedBookmarkButtonTagLeft�TopIWidthSHeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSharedBookmarkMoveToButtonTagLeft�TopiWidthSHeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick  TButtonUpSharedBookmarkButtonTag�Left�Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakTopakRight Caption   &Genväg...TabOrderOnClickShortCutBookmarkButtonClick    THistoryComboBoxLocalDirectoryEditLeft.TopWidth�HeightAnchorsakLeftakTopakRight DropDownCountTabOrder TextLocalDirectoryEditOnChangeDirectoryEditChangeSaveOn   THistoryComboBoxRemoteDirectoryEditLeft.TopIWidth�HeightAnchorsakLeftakTopakRight DropDownCount	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeDirectoryEditChangeSaveOn   TButtonLocalDirectoryBrowseButtonLeft�TopWidthKHeightAnchorsakTopakRight Caption   Blädd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop�WidthaHeightAnchorsakRightakBottom Caption   &Bokmärken...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPngImageListBookmarkImageList	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�����ɈEn?�m�&w�ܟG�@�3�xj�JK�b�P�����R?~�Ƹ�Y.DP�g���&��[�3�{�9����ƙ|����x$��~���p��i?	2nj��l�#$ƅb��W���f�|������.��l`����2 `���G��_W�_cp4���a�.����)�,��� lܾa�o��,V3c�SW�
�o�wɀ�T��ב��#(�[�a�U�f`g����)$2#~�Gр� ���l�Ԁ�@8uɀT/�?��l1�\`{��FJ���b��W�H�f`��I�+�.p8�`#"�����o�va���ÿ�X��?ܜ�Q�l%��	����a۝|R�Qm�b��)V���޽g0f���)܀O�4�7��2\����P�����O�ID  �/����>���I����ß?$�H)2��1|�r��~�d  m��7_��    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  iIDATx�c���?%�����ɈEn?�m�&w�ܟG�@�x��,"(ɿ�:� E���^|�y���Z�Z��h	I�H�{����+���yd3�k�6I�޽�*� F��	�$�y�y4�t.�|����;#��A��c�K�L�����3l�6@�L���Wms�?o����B#���G��0\:tw� Q	}5Q����©	�>����ǟ����13�j103~��-L!���20�X}�ǿ���HJr2���m�UȀd 
��~��p���~5=��9�0��)!�3��G�u���W3}k�`��,�(&BR�10|g��Oƣ��;F�s#�  6|�j���    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�c���?%�����ɈEn?�m�&w�ܟG�@��4�,f��,"(����GE��-�޽��W�x#^6��]��P��BQ���7��;�aw6�1���0���Ȓ���[3�V?d�@N��[y�$͛�M��Ne`�}9��J h���9'�Ȍ``�u�t�7�?�f@�ß���ۼ�2�����I�+��`�T����\�Q} ;t�%�>��N�j��e�>i^R��?��/~Տ�z)΍�  Tؚ�hƕ2    IEND�B`�  Left`Top� Bitmap
      TPngImageListBookmarkImageList120HeightWidth	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  KIDATx�c���?5#���D��0orMR��0�������IBc9 �o��d� ��w� �㋧�2���n�^�6F�RFF��� �:���O1�V�3r��Jf���;u��ѥ�/��3�
0�K��ad���×�_�<~��qS���D{���ّ��O1��81�����ׯ�� 6���9�����@6�؆;!�V�!��Ūf��lHnܶb�W��owC��cЌX��YLap��c`cc��i�a����K~|ޏ����(Z�bpP�B5��	���3~~9��%�赖�T�Xn>~b�{n7��og0\�ς5V��d�����r�����??��:d�j�5�rl,�^�1�>8��קh0��o=�`'"4�a��;�H��d����F���gXn��`�#����o�� ö{!Z{3����f`Dbo	��`�)�p������BL�a��gPf�559A�r�.��,�~f����=sA���? K���@uV$P������׊���C?Z�X����Td�Y��[�3��|���1$�x� }��%6 �$,a-)    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  /IDATx�c���?5#�����6��Hrk�y����$A�123�W��WՂ
�c�y`���׷~��(�C7�ʿдsW�r�C1���0��}������<N��w����$����f@a�(�����N�[h�.����͂C��c3�e �3�\��@��fA���f��mç�o(�����L��o�����C�_�e�mK�2���;{�F,f�٧��:���)�����~�v������o?ë�w��D�3Y���>y"ß����f�>(s^���o�����s6fxp�-��O<���W��i��Wg�8 �G���*�<"z����~�ƞ\��wN_cxp�N���^��*��8�tl�~?e���'���=�#�WN�c��擦oó�;{���2��V ��E�p�����a�)�j����]���U��������5�b�Hy��Í�Ϧ����"��&4��OL��P����/������}k���Y�#�)��ȹ?����%6 �L#�ēn\    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  [IDATx�c���?5#���D��0orMR��0�������!C��1�倬�����\�ީ�/�����!CQ��*wFN��X��C�S�]�@ȁG|��"l���hOv���h #���G`�[y�l�6��`�U�����ݰ Ơ�����s�`�Y���������kFY�o�bL=�g0��r�K����o�JL�s�~;��2b,�;o�j���B��^�Y�g�vL��~}��f ���w_�)y���~Bp|�!ķO��4��Ә�ߟ�53b����{X\�]�� 8�?��O��j����@)+2Фc>����A_b �$��l���    IEND�B`�  Left`Top� Bitmap
      TPngImageListBookmarkImageList144HeightWidth	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���_HSQ��q۝#��0�R�O�����Π?�$(��#�"D�7#������%��a�Ϳ��V�)��Q�`&����6w;��<�n�|�p�r~�����^"�"ֲ�� ��Q�%MT*Zi(��"�༵�j���h����T��ʿ]� ���b�3���nߗ༶�&Wve�����[��#�]���������Tޥ�nHݔ��Ή,��~�O�(s	���d���J�K&6�-��&��P�ղ1v�e.7Y �u��ӧ���C�(��ښ��Y�rbg�ڋ�|p1�g-�,�pvZ�k�q0��J���E�\Hx��GQ�����>8v��I[�Y��fcv�em����A8Zن�){�D1�4�0��@����!8R� �t�}7� =�R4����#̹;�}X���t
(���,p��]��H��	��i�r�e�8��~I��۴ �`V��	��c�C�W�}\�@��f3�aR��KJ�m�,Pt�~�p�ǯ7���I�D��@ �#-zeۧ�%���M���U�m�9�a���|��Fbf�I���>3�fkBAϊ	���,}��X(ao
*����t���kz�b���(�Ͻ�=�9�3>�Q�Z�FK-�@7ݲ%�Y�{Cǘ�`	�tg|�j���H���Cr�4�@�H	�:�w�m˄�1�fñ*����/�2Cen�`�� �«��?z    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
<  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-�з Dlj��f`b�d*�ɯ���QTX�/�- ��̸_��CT\U*��o���������<
"��M��/4�\��U5��a������=/n� ���s�j��-�5Q��Ex<����Ӡ0�-���;�Sk�\Z�W��O�eT�x,��]������m���**���_g�m`���9A�=����
�@��Ud8û'O>��`�qm����?�f�;5r���`�;��2Hh�2H�1���T|��?n�<�����Z����a0�of`b~����+���/~�6�w/^�-P�o��ph�&����>���_��gd@/����2\�����_���X0ܻ���$ ����8��X�|~����ݗ��Ih��9e&6y]�??�p-�� �]����S|k�-��gP0�b�ef���-i�Gc�si�Y����G��=Y� �֑L���?�'ϒ�+��oóG�;z�����1���1��r�Fl|�b~�e8}����G�`m�V�/��Ϡe ��o!l���wNm\����q ؂�
���E8����H��'>0<���Ŀ�q/X��V�������"���?v��3������lj�}���(�@-����+�*��_� %)c�^c�    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
9  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-�𰀑��as�����@!T%��0�������)��`K�4�p���f�Jf(
�:���⩫��8�b	���������f	)8�[��aA���������+�0�X��K5���i�L�|+�P����&���b��v5T�4�#��sfaZ�]������8°�?n��s`Z�U������d�S~�ܥ�x.b��i�>��{߼՘x�Oe���V���2�w�F,�3��v
�&�|��ў��0-pϪ`���2\#���gٞ�{0-�e���:C��#Ďﾁ%�u0�����A�Y�}j7�֞F��|�k #W#�=��>�d�]�W����l�6	Ղ-��G�RVT@���T?��[@K@s 	�E�35�    IEND�B`�  Left`TopBitmap
      TPngImageListBookmarkImageList192Height Width 	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
   �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  wIDATx���kHSa����L��X��ZT���Ce��)%i��
�[_*�~�@H���EW�2Z�ԩ�4�Nd����dB�[��]N�í�y�M�����{�=��}�ecA�p���`���H�'�D�C�ݚ�� |8�7 TI,N�X�'Y�����N���KE�}=�_�3�"�^RTѧ���}o���V�} PY�����|����QFDR��_xf�����ss�^H�F�-��1�c��Hu& �w�f��G{Gk��6> �>��jڂ��q'�;����x�p���':Mv�R��9F3�-V&0^�Z�"��׵W0?MC ,���tK�\93l ��1��J+��m�֝D��.d�! VI=_u�����y� ���"3y�4���d_=?��҄AW�G&��Y%P����[G�9�&L?9��'��@&�T��f1`��
����n�z��4��	`t@M�[1���*8������y�c�	@N��H�(g�'1�����R�S�+�j[�����o0��� ڋЩFJ꾵Q [K�;��c��MẶZyX��
���Al)������0B�a%�:�Ā�M���ބ��7A:Ǩ+�����58��m�8?i��0ꪐn�Jn���~-�|+�p��~MW;p�>7�\�6�Cj�����&hL ����T�D�{>S�������<4T٬"�Yy�ǃV�1N���� m�Tp�*��yw��}p��/�^d������1�!Cy2� ���!�[�8�w�lv1R��\.��X�I�g�t���VAǲLY�H���St�!��XS�Y��ێu�+������0w�`�Z]#@Hp���m�տ^ D��V7��|�զ �3��M*7ߠ*�    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  oIDATx��YLQ��QY�P1*Z4JDq�Ke	�.DB>�+�AM41�d���B�7L4j4��1FISæDD@ B��UKC-Pʴ�-�8�s[����M&s�̽�|�9��p�σ�>�*B�r��2�NaO����P�ax|q��čN'��`Nn�����[�5Z�̘<�0/9j��Ju�."Z��<�D̓���?5zL����̬��\����1�XE��@%f�QAG�͇�hMT�)����
Pr�:4@�~UX��1�ؾ;b�~k`1�a�!�����3��axePb�ɲ��<)Nu�팢 6��Y9X�2�"������C��!���]��������<.�!'BMl�憹�Ct�1�IL��@��b��p���Y~�O������RQw3G�R 2<hi䐰�� uQ'WH����`}������|Hs��M����@��kd�'x�}���4�Ȼ�lfI[������:W��P jR���I�|�:\�rO��O��c
�"Y&���+�7�i���F,]����b��=��Zf�~��w��9P����$o\
@�a��t$��@��ʬ���"K9����nE���F��Đ�S��!6^	�`	�0t���7=�h�����Wd �Hkw�bJ?Y�`�a�g��I�����Y�35��2�	�)����s�k����7�����p��cЭ�Ud�L���U�� vIT@�NbS_E����K��.nT��3�����K,X�
�6f�N@z�?��ͣ\��)9�L���qPΌ���%JA�LpTVm���s���f�y��|�	�^���s�R�ǿ˚[o0��ړ��3?��/�����w�Ǭ�E�v��� ? +L~?�
�    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?�@�Q�: � FFF��",r{�α¡�ȏ?���~�k6����E�[�>�D�*���G'0�8��ͯ�q5���Y֜���ih*#+'VͿ|c8�z�߿_���6<;GUln�����#���׀���0\ݷ�� 8�[�����;'�k0Q`��@0�t�}�Mpp�%����P����ghj��v��.�����&$��Te�3��J�3|}��h�It��9s�;��x=���;H���Ca�܅��Y������8!5D0���]B��~|ޏ�@�����+�;�#:ï/�������yk	8 �����$?���H�9�����Jpc���y��;�=���Ϗ�DY���ՠ����E�yަ��q9`~��'3����aB����=�~��:��v�ϧĉ�}�@I�[�����&V�����`�	t�oTI*Y�v? Pfi�R��l�6	��>�<4@{���<��ꀁ�  Iӯ�v �	    IEND�B`�  Left`Top@Bitmap
       TPF0TLoginDialogLoginDialogLeft_Top� HelpType	htKeywordHelpKeywordui_loginBorderIconsbiSystemMenu
biMinimizebiHelp Caption
InloggningClientHeight�ClientWidthiColor	clBtnFaceConstraints.MinHeight�Constraints.MinWidthX
ParentFont	
KeyPreview	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShowPixelsPerInch`
TextHeight TPanel	MainPanelLeft Top WidthiHeightiAlignalRight
BevelOuterbvNoneTabOrder  TPanelContentsPanelLeft Top WidthiHeight@AlignalClient
BevelOuterbvNoneTabOrder Visible
DesignSizei@  	TGroupBoxContentsGroupBoxLeftTopWidth[Height1AnchorsakLeftakTopakBottom CaptionContentsGroupBoxTabOrder 
DesignSize[1  TLabelContentsLabelLeftTopWidthHeightCaptionNamn:ShowAccelChar  TEditContentsNameEditLeftBTopWidthHeightAnchorsakLeftakTopakRight TabOrder TextContentsNameEdit  TMemoContentsMemoLeftTop*WidthDHeight� AnchorsakLeftakTopakRightakBottom Lines.StringsContentsMemo TabOrder    TPanel	SitePanelLeft Top WidthiHeight@AlignalClientAnchorsakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSizei@  	TGroupBox
BasicGroupLeftTopWidth[Height� AnchorsakLeftakTopakRight CaptionSessionTabOrder 
DesignSize[�   TLabelLabel1LeftTopHWidth7HeightCaption   &Värdnamn:FocusControlHostNameEdit  TLabelLabel2Left� TopHWidth?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlPortNumberEdit  TLabelUserNameLabelLeftTopzWidth7HeightCaption   &Användarnamn:FocusControlUserNameEdit  TLabelPasswordLabelLeft� TopzWidth2HeightCaption   &Lösenord:FocusControlPasswordEdit  TLabelLabel22LeftTopWidth>HeightCaption&Filprotokoll:FocusControlTransferProtocolCombo  TLabel	FtpsLabelLeft� TopWidth7HeightCaption&Kryptering:FocusControl	FtpsCombo  TLabelWebDavsLabelLeft� TopWidth7HeightCaption&Kryptering:FocusControlWebDavsCombo  TEditEncryptionViewLeft� Top'Width� HeightTabOrderOnChangeTransferProtocolComboChange  TEditTransferProtocolViewLeftTop'Width� HeightTabOrderOnChangeTransferProtocolComboChange  TEditHostNameEditLeftTopYWidth� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderTextHostNameEditOnChange
DataChangeOnExitHostNameEditExit  TEditUserNameEditLeftTop� Width� Height	MaxLength� TabOrderTextUserNameEditOnChange
DataChange  TPasswordEditPasswordEditLeft� Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextPasswordEditOnChange
DataChange  TUpDownEditPortNumberEditLeft� TopYWidthRHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChangePortNumberEditChange  	TComboBoxTransferProtocolComboLeftTop'Width� HeightStylecsDropDownListTabOrder OnChangeTransferProtocolComboChangeItems.StringsSFTPSCPFTPWebDAV	Amazon S3   	TComboBox	FtpsComboLeft� Top'Width� HeightStylecsDropDownListTabOrderOnChangeTransferProtocolComboChangeItems.StringsIngen krypteringTLS/SSL Implicit encryptionXTLS/SSL Explicit encryptionX   	TComboBoxWebDavsComboLeft� Top'Width� HeightStylecsDropDownListTabOrderOnChangeTransferProtocolComboChangeItems.StringsNo encryptionXTLS/SSL Implicit encryptionX   TPanelBasicFtpPanelLeftTop� WidthDHeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder	 	TCheckBoxAnonymousLoginCheckLeft Top Width� HeightCaption&Anonym inloggningTabOrder OnClickAnonymousLoginCheckClick   TPanelBasicSshPanelLeftTop� Width[Height AnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
  TButtonAdvancedButtonLeft� Top� WidthbHeightActionSessionAdvancedActionAnchorsakRightakBottom StylebsSplitButtonTabOrderOnDropDownClickAdvancedButtonDropDownClick  TButton
SaveButtonLeftTop� WidthbHeightActionSaveSessionActionAnchorsakLeftakBottom StylebsSplitButtonTabOrderOnDropDownClickSaveButtonDropDownClick  TButtonEditCancelButtonLefttTop� WidthRHeightActionEditCancelActionAnchorsakLeftakBottom TabOrderOnDropDownClickSaveButtonDropDownClick  TButton
EditButtonLeftTop� WidthbHeightActionEditSessionActionAnchorsakLeftakBottom TabOrderOnDropDownClickSaveButtonDropDownClick   	TGroupBox	NoteGroupLeftTop� Width[HeightFAnchorsakLeftakTopakRightakBottom Caption
AnteckningTabOrder
DesignSize[F  TMemoNoteMemoLeftTopWidthMHeight.TabStopAnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneLines.StringsNoteMemo 
ScrollBars
ssVerticalTabOrder     TPanelButtonPanelLeft Top@WidthiHeight)AlignalBottom
BevelOuterbvNoneTabOrderOnMouseDownPanelMouseDown
DesignSizei)  TButtonLoginButtonLeftKTop
WidthbHeightActionLoginActionAnchorsakRightakBottom Default	ImagesActionImageListModalResultStylebsSplitButtonTabOrder OnDropDownClickLoginButtonDropDownClick  TButtonCloseButtonLeft� Top
WidthRHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  TButton
HelpButtonLeftTop
WidthRHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPanel
SitesPanelLeft Top Width HeightiAlignalClient
BevelOuterbvNoneTabOrder
DesignSize i  	TTreeViewSessionTreeLeftTopWidth�Height8AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesSessionImageListIndentParentDoubleBufferedParentShowHint	RowSelect	ShowHint	ShowRootSortTypestBothTabOrder OnChangeSessionTreeChange
OnChangingSessionTreeChangingOnCollapsedSessionTreeExpandedCollapsed	OnCompareSessionTreeCompareOnContextPopupSessionTreeContextPopupOnCustomDrawItemSessionTreeCustomDrawItem
OnDblClickSessionTreeDblClick
OnDragDropSessionTreeDragDropOnEditedSessionTreeEdited	OnEditingSessionTreeEditing	OnEndDragSessionTreeEndDragOnExitSessionTreeExitOnExpandingSessionTreeExpanding
OnExpandedSessionTreeExpandedCollapsed	OnKeyDownSessionTreeKeyDown
OnKeyPressSessionTreeKeyPressOnMouseDownSessionTreeMouseDownOnMouseMoveSessionTreeMouseMoveOnStartDragSessionTreeStartDrag  TStaticTextSitesIncrementalSearchLabelLeftTop0Width�HeightAnchorsakLeftakRightakBottom BorderStyle	sbsSingleCaptionSitesIncrementalSearchLabelShowAccelCharTabOrderVisible  TButtonManageButtonLeft�TopJWidthbHeightAnchorsakRightakBottom Caption&HanteraTabOrderOnClickManageButtonClick  TButtonToolsMenuButtonLeftTopJWidthbHeightAnchorsakLeftakBottom Caption&VerktygTabOrderOnClickToolsMenuButtonClick   TPanelShowAgainPanelLeft TopiWidthiHeightAlignalBottom
BevelOuterbvNoneTabOrderOnMouseDownPanelMouseDown
DesignSizei  	TCheckBoxShowAgainCheckLeftTop WidthQHeightAnchorsakLeftakTopakRight CaptionO   &Visa inloggningsdialogrutan vid start och när den sista sessionen är stängdChecked	State	cbCheckedTabOrder    TActionList
ActionListImagesActionImageListOnUpdateActionListUpdateLeft,Top TActionEditSessionActionCategorySessionsCaption	&Redigera	OnExecuteEditSessionActionExecute  TActionSaveAsSessionActionCategorySessionsCaption
&Spara somShortCutA�  	OnExecuteSaveAsSessionActionExecute  TActionSaveSessionActionCategorySessionsCaption	&Spara...	OnExecuteSaveSessionActionExecute  TActionDeleteSessionActionCategorySessionsCaptionTa &bort...
ImageIndex	OnExecuteDeleteSessionActionExecute  TActionImportSessionsActionCategorySessionsCaption&Importera...	OnExecuteImportSessionsActionExecute  TActionLoginActionCategorySessionCaptionLogga in
ImageIndex 	OnExecuteLoginActionExecute  TActionAboutActionCategoryOtherCaption&Om...	OnExecuteAboutActionExecute  TActionCleanUpActionCategoryOtherCaption&Rensa applikationsdata...	OnExecuteCleanUpActionExecute  TActionResetNewSessionActionCategorySessionsCaption   Å&terställ	OnExecuteResetNewSessionActionExecute  TActionSetDefaultSessionActionCategorySessionsCaption   Sä&tt som standard	OnExecuteSetDefaultSessionActionExecute  TActionDesktopIconActionCategorySessionsCaptionSkrivbords&ikon	OnExecuteDesktopIconActionExecute  TActionSendToHookActionCategorySessionsCaption"   Utforskarens 'Skicka till'-genväg	OnExecuteSendToHookActionExecute  TActionCheckForUpdatesActionTagCategoryOtherCaption   Sök efter &uppdateringar
ImageIndex?	OnExecuteCheckForUpdatesActionExecute  TActionRenameSessionActionCategorySessionsCaption	Byt &namn
ImageIndex	OnExecuteRenameSessionActionExecute  TActionNewSessionFolderActionCategorySessionsCaptionN&y katalog...
ImageIndex	OnExecuteNewSessionFolderActionExecute  TActionRunPageantActionCategoryOtherCaption   Kör &Pageant	OnExecuteRunPageantActionExecute  TActionRunPuttygenActionCategoryOtherCaption   Kör PuTTY&gen	OnExecuteRunPuttygenActionExecute  TActionImportActionCategoryOtherCaption'   Importera/Återställ &konfiguration...	OnExecuteImportActionExecute  TActionExportActionCategoryOtherCaption-   &Exportera/Säkerhetskopiera konfiguration...	OnExecuteExportActionExecute  TActionPreferencesActionCategoryOtherCaption   &Inställningar...	OnExecutePreferencesActionExecute  TActionEditCancelActionCategorySessionCaption&Avbryt	OnExecuteEditCancelActionExecute  TActionSessionAdvancedActionCategorySessionCaption&Avancerad...	OnExecuteSessionAdvancedActionExecute  TActionPreferencesLoggingActionCategoryOtherCaption&Loggning...	OnExecutePreferencesLoggingActionExecute  TActionCloneToNewSiteActionCategorySessionCaption&Klona till ny webbplats	OnExecuteCloneToNewSiteActionExecute  TActionPuttyActionCategorySessionCaption   Öppna i &PuTTY
ImageIndexSecondaryShortCuts.StringsShift+Ctrl+P ShortCutP@	OnExecutePuttyActionExecute  TActionPasteUrlActionCategorySessionsCaptionKlistra in sessions-&URLShortCutV@	OnExecutePasteUrlActionExecute  TActionGenerateUrlAction2CategorySessionsCaption&Skapa sessions-URL/kod...	OnExecuteGenerateUrlAction2Execute  TActionCopyParamRuleActionCategorySessionsCaption#   Överföringsinställnings&regel...	OnExecuteCopyParamRuleActionExecute  TActionSearchSiteNameStartOnlyActionCategoryOtherCaption$   Endast &början av webbplatsens namn	OnExecute$SearchSiteNameStartOnlyActionExecute  TActionSearchSiteNameActionCategoryOtherCaption&Varje del av webbplatsens namn	OnExecuteSearchSiteNameActionExecute  TActionSearchSiteActionCategoryOtherCaption   Alla &fält för webbplatsen	OnExecuteSearchSiteActionExecute  TActionSessionRawActionCategorySessionCaption   Redigera Raw-inställningar...	OnExecuteSessionAdvancedActionExecute   
TPopupMenuToolsPopupMenuLeft� TopM 	TMenuItemImport1ActionImportSessionsAction  	TMenuItemN3Caption-  	TMenuItemImportConfiguration1ActionImportAction  	TMenuItemExportConfiguration1ActionExportAction  	TMenuItemCleanup1ActionCleanUpAction  	TMenuItemN2Caption-  	TMenuItemPageant1ActionRunPageantAction  	TMenuItem	Puttygen1ActionRunPuttygenAction  	TMenuItemN1Caption-  	TMenuItemCheckForUpdates1ActionCheckForUpdatesAction  	TMenuItemN4Caption-  	TMenuItemPreferences1ActionPreferencesAction  	TMenuItemAbout1ActionAboutAction   TPngImageListSessionImageList	PngImages
BackgroundclWhiteNameUnusedPngImage.Data
b   �PNG

   IHDR         ��h6   tRNS �   ���/�   IDATx�c����8�aT���  �E�/UY"    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
J  �PNG

   IHDR         ��h6   tRNS � � �7X}   �IDATx�c���?)��d�IϞ�$�NJR|�� ��ދ������������P�?�rA��S�@5L��谿���p�.T��IC�� Q�:	R��d�1�:���5HHP��_�����������ן�����j���k�Ƽ��������T`z��(����������_(]���`���`����`�����C}d5jx|�TC`dʓg�I�i��d��gC�DOKp�J��6�S+ ����>�7    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  iIDATx�c���?%�����ɈEn?�m�&w�ܟG�@�x��,"(ɿ�:� E���^|�y���Z�Z��h	I�H�{����+���yd3�k�6I�޽�*� F��	�$�y�y4�t.�|����;#��A��c�K�L�����3l�6@�L���Wms�?o����B#���G��0\:tw� Q	}5Q����©	�>����ǟ����13�j103~��-L!���20�X}�ǿ���HJr2���m�UȀd 
��~��p���~5=��9�0��)!�3��G�u���W3}k�`��,�(&BR�10|g��Oƣ��;F�s#�  6|�j���    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�c���?%�����ɈEn?�m�&w�ܟG�@��4�,f��,"(����GE��-�޽��W�x#^6��]��P��BQ���7��;�aw6�1���0���Ȓ���[3�V?d�@N��[y�$͛�M��Ne`�}9��J h���9'�Ȍ``�u�t�7�?�f@�ß���ۼ�2�����I�+��`�T����\�Q} ;t�%�>��N�j��e�>i^R��?��/~Տ�z)΍�  Tؚ�hƕ2    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
/  �PNG

   IHDR         ��h6   tRNS � � �7X}   �IDATx�c���?)��d�A-���!F���ȥ�Ռ<f���h8�����~�������Ԁ�0oѪ��0	��Ahx~�Ͱ����m�%�J����t�P��J� �-K���ؠ	�9�B5��ӅfX����h�J.eP7wv�8u(�a�d ��UǊì���ˡ�l�@3l���y��h�:^P�7���M�p"3�M�з�!-ٟ�x�5w#NOcPO���HM� WՌ�\[    IEND�B`� 
BackgroundclWindowNameWorkspace closedPngImage.Data
b   �PNG

   IHDR         ��h6   tRNS �   ���/�   IDATx�c����8�aT���  �E�/UY"    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ���``d���)��!�WL�Lɟ?���͸�H����d��>����7Y��~��[��+����89�l��׷��fx����/�=xe��+�^��g�����3T�c���c�d����쵇N_�߸�+������P�"6ظ���M|����M8�X��g`�}������z�d��)��%�3 ���H��d��w>3�>w�!�ǂAJT��ś��w�e�q������OY���1�ç��Na�a`fbb��g�u��敝�~ W���_�5 �f`x��1ã�w�5~���p���?��Vv��(�^������>1����?÷_@��l�b�ѵ�^љvn@^����|���������3���=f.�f8}p+<���6lfx����M���$_L��� ���DLd5�6������D���ph�� l*@����m�qiD� :�lV�B    IEND�B`� 
BackgroundclWindowNameOpen new session closedPngImage.Data
r   �PNG

   IHDR         ��h6   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?)�qTè�� ��/�Ǭ�Y    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�   �PNG

   IHDR         ��h6   tRNS � � �@�   bIDATx�c�����H����g�_T'%)��pH���w��K54D��:<���d5jx|�TC`dʓg�	j@�4ZZ2+���!F��d�� Mɩ �ROqe�!�    IEND�B`�  Left,Top� Bitmap
      
TPopupMenuSaveDropDownMenuLeftTop 	TMenuItemSaveSessionMenuItemActionSaveSessionActionDefault	  	TMenuItemSaveAsSessionMenuItemActionSaveAsSessionAction  	TMenuItemN7Caption-  	TMenuItemSetdefaults1ActionSetDefaultSessionAction   
TPopupMenuManageSitePopupMenuImagesActionImageListLeft�Top 	TMenuItem
Shellicon1Caption	WebbplatsEnabledVisible  	TMenuItemSiteLoginMenuItemActionLoginActionDefault	  	TMenuItemOpeninPuTTY2ActionPuttyAction  	TMenuItemN10Caption-  	TMenuItemEdit1ActionEditSessionAction  	TMenuItemDelete1ActionDeleteSessionAction  	TMenuItemRename1ActionRenameSessionAction  	TMenuItemSiteClonetoNewSiteMenuItemActionCloneToNewSiteAction  	TMenuItemGenerateSessionURL1ActionGenerateUrlAction2  	TMenuItemN5Caption-  	TMenuItemSetdefaults2ActionSetDefaultSessionAction  	TMenuItemN6Caption-  	TMenuItem
Newfolder1ActionNewSessionFolderAction  	TMenuItem
Shellicon2CaptionIkon webbplatsEnabledVisible  	TMenuItemDesktopIcon2ActionDesktopIconAction  	TMenuItemExplorersSendToShortcut2ActionSendToHookAction  	TMenuItemOptions1Caption
AlternativEnabledVisible  	TMenuItemIncrementalSearch1Caption   Inkrementell sökning 	TMenuItemSearchSiteNameStartOnly1ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemSearchSiteName1ActionSearchSiteNameAction	RadioItem	  	TMenuItemSearchSite1ActionSearchSiteAction	RadioItem	    
TPopupMenuManageFolderPopupMenuImagesActionImageListLeft�TopM 	TMenuItem	MenuItem1CaptionWebbplatskatalogEnabledVisible  	TMenuItemLogin5ActionLoginActionDefault	  	TMenuItemN11Caption-  	TMenuItem	MenuItem3ActionDeleteSessionAction  	TMenuItem	MenuItem4ActionRenameSessionAction  	TMenuItem	MenuItem5Caption-  	TMenuItem	MenuItem6ActionNewSessionFolderAction  	TMenuItem	MenuItem7CaptionIkon webbplatskatalogEnabledVisible  	TMenuItem	MenuItem8ActionDesktopIconAction  	TMenuItemOptions3Caption
AlternativEnabledVisible  	TMenuItemIncrementalSearch3Caption   Inkrementell sökning 	TMenuItemBeginningofSiteNameOnly2ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemAnyPartofSiteName2ActionSearchSiteNameAction	RadioItem	  	TMenuItemAllMajorSiteFields2ActionSearchSiteAction	RadioItem	    
TPopupMenuManageNewSitePopupMenuImagesActionImageListLeft� Top�  	TMenuItem
MenuItem12CaptionNy webbplatsEnabledVisible  	TMenuItemLogin2ActionLoginActionDefault	  	TMenuItemOpeninPuTTY3ActionPuttyAction  	TMenuItemN8Caption-  	TMenuItem
MenuItem13ActionSaveAsSessionAction  	TMenuItemReset1ActionResetNewSessionAction  	TMenuItemPaste1ActionPasteUrlAction  	TMenuItemGenerateSessionURL2ActionGenerateUrlAction2  	TMenuItem
MenuItem21Caption-  	TMenuItem
MenuItem22ActionSetDefaultSessionAction  	TMenuItem
MenuItem16Caption-  	TMenuItem
MenuItem17ActionNewSessionFolderAction  	TMenuItemOptions2Caption
AlternativEnabledVisible  	TMenuItemIncrementalSearch2Caption   Inkrementell sökning 	TMenuItemBeginningofSiteNameOnly1ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemAnyPartofSiteName1ActionSearchSiteNameAction	RadioItem	  	TMenuItemAllMajorSiteFields1ActionSearchSiteAction	RadioItem	    
TPopupMenuManageWorkspacePopupMenuImagesActionImageListLeft�Top�  	TMenuItem	MenuItem2Caption	ArbetsytaEnabledVisible  	TMenuItemLogin3ActionLoginActionDefault	  	TMenuItemN9Caption-  	TMenuItem
MenuItem10ActionDeleteSessionAction  	TMenuItem
MenuItem11ActionRenameSessionAction  	TMenuItem
MenuItem18CaptionIkon arbetsytaEnabledVisible  	TMenuItem
MenuItem19ActionDesktopIconAction  	TMenuItemOptions4Caption
AlternativEnabledVisible  	TMenuItemIncrementalSearch4Caption   Inkrementell sökning 	TMenuItemBeginningofSiteNameOnly3ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemAnyPartofSiteName3ActionSearchSiteNameAction	RadioItem	  	TMenuItemAllMajorSiteFields3ActionSearchSiteAction	RadioItem	    
TPopupMenuSessionAdvancedPopupMenuLeft� Top 	TMenuItemSession1CaptionSessionEnabledVisible  	TMenuItem	MenuItem9ActionSessionAdvancedActionDefault	  	TMenuItemEditRawSettings1ActionSessionRawAction  	TMenuItemTransferSettingsRule1ActionCopyParamRuleAction  	TMenuItem
MenuItem14Caption   Globala inställningarEnabledVisible  	TMenuItemPreferencesLoggingAction1ActionPreferencesLoggingAction   TPngImageListActionImageList	PngImages
BackgroundclWindowNameLoginPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��o�d  �IDATx�cTh��!������ ���g*�|��oIavfR�3���������.�/�/\㰗A�S���ߟ0�p��]|� 6 ���1�[V[������⚂`��w,6����F=]������b �����CU �
��`�N�~��C����/�@V�������N=zL����a��.���3���,n�Z	,���G����"�����jO2�	<�`�\,���g�2<�c��gj�2�9�`�D,����|��.�?�{a�����炽 �_(����+� 1N���'��d��ǟ2��f����`d5_^}��%�����A{�4���8���H÷�_Q\���ۻ8����3�3hN���j~|�1���,�'���^�|z�������783��3�0222��������_pf�(; 1bҩCo��    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATxڅ�]HSa�g�meVt��6J�����.�0��""
��� �nv�]bA݈�1�>�"��8��bj�)i���)��R��<����ak{�����=���#��Qy`H��GP����XPAQ��G�M��.�%+�r��x�:"�Ǎ&/���;�����Of��7b���%n,%*���Dbs�����'(��c�f�>��,|��zMg��̀��2ŵ���1�������AL^�׵�D��lK�fY��3;��ؿ�$3�~���)Z'v�
?�)n���c�F��܀$�]���f&g��� O�-���������^!e��sa4ф���O��I�n����p[E�|���,TK�*/�*K�Ect>����(��k�W�F�cI��~�شX?
uW�����P�Z�f?O{c.������f](���̿��n���K��+<���'f���ׅ#�J�|�5����ʸ�� �"�Mg�)��01%�X���L6)WH������5�(�    IEND�B`� 
BackgroundclWindowNameRenamePngImage.Data
y  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ���+-+���ɋ�'>,`$Es������'�uT����p��`�Ḫ\���`����:?���G�h6����h������_��'6nk��v~+��^�w��Z����GW�}[� F�@C����"g��op�����������y�$G�痛�Է2P���5ÍK7�m�U����Qln�p
�Z�)`��������W?�
�g/���fF���&��l���y�p��%�E�QՀXؒ�ՀgW�2Hrng`�Nexz���U��A@�._3b���$���yF���?d �A��5-1v��^�aP�bH؀���`����06\Z�ɠ������YQ�(nQ@��L�I �,`��A`Ru:���&��e(��4�A���U�3�/d�U�c�|��5�1e-�|��X��l@gY1��w-���  �����i�    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
z  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�]HSaǟ�M�9�۔�t�ϴYJhe H!E7xQN*���Oꦫ��i	]TDA�`XMLYY:�3C��<�̹������$Q���}���<����B�'�� p��S!�nPO���V���|�J����=*I^��qN��^g�F˸ϯ,�m���wq'�Y���vǆ��	<C�vAr� �����RU�(.��b��y�D"��C����ss�4E�*/�;����y���/���7��YL��7WI HQx�i8�Jɻ	���Tߦ�{����&atb꣬��:67U	���\���﨩��`^����H��k+J,vk>��g�;��f�$�T��"^ m<{���9�XUM������d��0�O�irE"���V �����Z���3�lO��O�H ���X6w ��Ȼ��6ڨשg��2��7eF_���'t4yc���dqw!���͌Z�G�,^��`0�
p�gϲ4}��X�E\�e���4Bɭ�3�x�&S�X�Q��H.�F�*GQgx��8�AT�
j�m|����c��+��L>������5�|�^o2�TbK���S.Q���m$���i-6���Lɝح �V
��:�fF�i�\���VX�`(�~]I�v�4 �a�D�X�V,�}�{�%J���L]&}������T��Zp�7����x �D����LB����k�RFfP    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ���bd`���z�����/�j���?,|���o2c@X٬Yq����|<�����,,L�~��Zѝ������d�"���Mߑs�_�0�����n}>n�w�1�x������+�2�0nn���Ym�������&�d�72Ԑg���e�d���;ì��N_{X��+��qS��Uk%-!1.޽�ưi���B,̬��M�YY��g`�q�
�������d�WY���A�a��$�XosIQ��?0��}������1�_6 _ ~�+�p���AD������AB������=m�� �[y�G/<a8t����
��o?l� �wCu�R$�S~_G�����Rw^�2�x�!��8����cՀC�y�Y��GH�z10�y���?��P�͋.��h����#�dW`q����9+00���%��� *v��KT|R�1���c˜9(|Ҽ$������<�a���?)z1  �O�ہZ�    IEND�B`�  Left)Top� Bitmap
      
TPopupMenuLoginDropDownMenuImagesActionImageListLeftTopM 	TMenuItemLogin1ActionLoginActionDefault	  	TMenuItemOpeninPuTTY1ActionPuttyAction   TPngImageListSessionImageList120HeightWidth	PngImages
BackgroundclWindowNameUnusedPngImage.Data
v   �PNG

   IHDR         �Z   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?��qT��Qͣ�V3 O�;ه>�    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��o�d  rIDATx�cd�2`������g��1�f�=}p�	����]�����1����J�G���`�@<�6�h #���v��PEh��������O?�3l�F50�m=�uh.�����l �	��2/������Aٟ���}����;��0Tpi.��6 �� ��W��_�3����dpav��q`������ￄ��s��"%�~��/?30|�I�A0pzF ��~囀��醁�����Zfo"� 8>��@���xt�/��Ύ�$r�v.��:�̰w�~��&v�'�,3J\L����jN���QTG��'�o�ՃU���"����S9aqi�>ЋJ��������3�]��BJ  3 �{W�_    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  /IDATx�c���?5#�����6��Hrk�y����$A�123�W��WՂ
�c�y`���׷~��(�C7�ʿдsW�r�C1���0��}������<N��w����$����f@a�(�����N�[h�.����͂C��c3�e �3�\��@��fA���f��mç�o(�����L��o�����C�_�e�mK�2���;{�F,f�٧��:���)�����~�v������o?ë�w��D�3Y���>y"ß����f�>(s^���o�����s6fxp�-��O<���W��i��Wg�8 �G���*�<"z����~�ƞ\��wN_cxp�N���^��*��8�tl�~?e���'���=�#�WN�c��擦oó�;{���2��V ��E�p�����a�)�j����]���U��������5�b�Hy��Í�Ϧ����"��&4��OL��P����/������}k���Y�#�)��ȹ?����%6 �L#�ēn\    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  [IDATx�c���?5#���D��0orMR��0�������!C��1�倬�����\�ީ�/�����!CQ��*wFN��X��C�S�]�@ȁG|��"l���hOv���h #���G`�[y�l�6��`�U�����ݰ Ơ�����s�`�Y���������kFY�o�bL=�g0��r�K����o�JL�s�~;��2b,�;o�j���B��^�Y�g�vL��~}��f ���w_�)y���~Bp|�!ķO��4��Ә�ߟ�53b����{X\�]�� 8�?��O��j����@)+2Фc>����A_b �$��l���    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
S  �PNG

   IHDR         ��   	pHYs  �  ��o�d  IDATx�cd�2`�����02�צ�i�.3*Į���D�Vm�� 6PHL�*�{�b��rG���E�����
H�w����Q��Zɛ ^���p���V���@j@@/m3���3|��BÌ-OO����m0�c�����Ԁ�i��S���B����L��<uL���`e� 5 `��b��~O��оp;�������������q�0]5pW�U\�V�b`�� U\w���m��T1Ы|'�C�� ������	�    IEND�B`� 
BackgroundclWindowNameWorkspace closedPngImage.Data
v   �PNG

   IHDR         �Z   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?��qT��Qͣ�V3 O�;ه>�    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��o�d  kIDATxڥ�_HSQǿw�n�%�?�ʌ����A�dd�^��*��$z�(zQ���$\a�=�l�G�M3tS��hF�ess�m�������֘��\���������ˡ�54��(M��X��k��9j-��w����h��w��b���4��3�{@<���?D�H�q�P�֣���RZ�LؠT��%���%��������+���B��v��M�Ր24�*v@H��dR�����ׯM[ǁqh�O�?�-�U����Z�#1Pd5�H�os���^���$��ݘJ�O�xa�ŨՈ�{�(R����L�<h�6�e���{���}p�����kbڊ�W�qʢB�O�0=3�?�~�c:	���'�FG��<!���h��+����A��[�~;oD��s�b��$�R�;"(@��b,�_R,�\$�P�Џ>T�u�Q��ƞ���9UæV95
l8�M�y?�̐��bK%l�3�@�]��*�<,���Ng���J��S}&�ȍ޼�;OeOj���}!�5W�g���ju���'!�_G�Vs���M��<�~N9r��:IJ0I���ȥ��M��%���Ε�����{ok��9����/>6��'M�    IEND�B`� 
BackgroundclWindowNameOpen new session closedPngImage.Data
v   �PNG

   IHDR         �Z   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?��qT��Qͣ�V3 O�;ه>�    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�   �PNG

   IHDR         ��   	pHYs  �  ��o�d   �IDATx�cd�2`������g��1�f�=}p�	����n��43{�����8�tvt$ِc�s����d����#4��>	d�Q����N�9�՜`i#�������M�z�J���R�߾|�"',.c�zQ�X�[9���}��aF�� �]H	  �Stj     IEND�B`�  Left� Top� Bitmap
      TPngImageListActionImageList120HeightWidth	PngImages
BackgroundclWindowNameLoginPngImage.Data
/  �PNG

   IHDR         �Z   tRNS �  $�ݺ:  �IDATx�c|+��@.`j^�*k���~����=Ϻ4"lH�U�W~U.6.V"5������o�&r�4g��6�˭��+�)�U���OB:O/�9;U�YRW���-��jX5å�_~��,�%Wq���&U���R/��Ch���8p�|�J��Ԏ5~�G��2^�x��,�* Wq:���Ze �����s5���@�2�����,�ć��3a�!�}Ov������=D�d�"����'�fAy�s�p�Pg�骽���-W ����Y@��|�C<�[NV�}���p�<H���f>In4�A{no>Q���{���B9 ����<b\pm���Γ�@��V�~�M
����B3�\ŕ��:s��]f7)����s R@��7?�9��*��?Ӛ)���p���"4s��U\�z�9M�f�ԏO��ٸYjo�)>9���|z������7T30K�e�����@���?�?h���0 R&  �C��N��    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
Y  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڕ�mHSQ���9��d�8��|[*���C���0�
��B��>�("
��@0A?d$����/���niM͖/9M͖��ܽ�{�a]7����������\��������H ɽ�rp��#|�s# �0Z����?I���G�Q r�"X���u a�u�`�o�\ʖ^.��p?�!�ʅ�C�R�iw<I�$ �C��J�nU���Ba�ź ������C�1���I���<�0�`�i����KD��ݰY�0��P����� su��?�H
�+f1��I�B��'�03�^ƣ���!���VE����
e�=��FIu��$�T��mDf�;�	e���;�x�ZF�(��dؼ� E�fYhy�_�D�~{4ڧ�E�Q��=�6�}.�c�I�Y��#��j�2?�_���
m�j��V^��xx���g�q�ii�����Ƈ�W_��a%��j|��d��^c�K�o�."�X��尽��`[^�o@�`������&�կ3�Ad�Z0b@{�u4V�� ^'<{����3��l�YH1�� �p�#�� ��$0�X�w��&TL��Fe�.'&��0��`Q��5I��s�"1�v!����ɀE{����&	�J��e��y�-�=�I��'��Wz���Y`V�_�� �mcN�ڻ�    IEND�B`� 
BackgroundclWindowNameRenamePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��o�d  �IDATxڝ�]H�Q���s-M-Ԗ.%��XI��d�$ˌʋ(?iX�D&�EZT䠰ش	tم*�b���:��iKc��̡��� j6���{�s��wq�˂�� v8�+w~�&��;����|[y<q��/��
�JCO��Dv��'0�Dup�yt�l'S&��蛵4UX�W}��.ʎ�Db���ptu�-A5`�|vm۞��DՄ%ݱ�%���`|��jy�R��R��a;�i���� tZ�z��ޓɎ;���;��̓9���6,��a�<u߯݅�Ġ�g���'���3����ߣ���*�����[3��9�-�ԁR��͘7��^m��&�����5H"��^UĎ$���w��wO��������<�.mFAzg�>����O�zg��γ������c8��-��~�3��U�
��d��b��~TJ�nl�0�-F��L���i���d��6��/�(V@E��zR�P��@�$ýX�V����u���W#&�1��݂�`��TS(���Z�h���o����/.a�E�^�g��u�L����5�k�y٩0��
�B���^$��")a
U҇p�IN�@��5�����`��Vm1.5+���#� {���J�_n /(�#FB�^sfM�r�F������1������    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
R  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڭ�[lU��̙���em;n]ZiI@
mll-]�Q�$�DbBB⛁��㛉>ߌ)-}�1F�O�Ub��K�\KK�.�ݖ]螹�\<3kW[���y�9g�{��7��s� D�7�0��ܼ�����^>$�	�ל�z$���`kd�_��-��Q_�s�j�p4��Ǖ��b�!d[��!�B!�(��R�.8~���w9BvP�Y�HR;��/���JKKd2�`>_��!!x8&�ŎnM=���{�<}���(���^u�r��g��;��5��ޜ�3�nڮ׳O�n��$=ųxlK�f1W�=��vz�wJ��QՃ�6c�vs_�t��q��������ߧ�S�2�.����M땵�x����g'a�����?a���'7qu1�,�L\�,�y1�������`�5�q?��<�v}c"����M����ɶ�H�@tF'�˶�үiǗ��V���?��X{kS5�J��<�i����t��}�|��b�QY~k����п׭���9����OWVU�V�ڨN���ln�0���a�Y������/�b<žn��vѶ`��U�&�4��\�X��
*���! ���c���lm�`>X?�P���
��S��B�����}�y�`%7dm��1��];{�s�����2��I����Rtr�4���5mn8 ��<�?o"����)U��eϕ���wM��(f>J�>�`3��4}J#�ַ�Up��`=�>�������j��G�$K�C��f�nh�( ���Mf����a!��<��Ž9�9\.�i��=��^Y�!I��#����������>-:n}�p5�JA��A�ߛ�/�_�o�v|��6��7M#κ�Sv��3���T�r�v���x��F{��w����X��>��6w�����    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
2  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ��6�1*J�2��J�F�c$����^�
�[����p��˨?��cffQ{���a�-�bb�i:��5J
��V�a����A��������ջ/�`77H��ga�t�	�g����mx��)����ͱ3�˜�����PC���߿`��X�J��0<}�ޑb�Y}3m%3�q�/�d�w��U�? �60��J��2PN�g���#�9 ��ɰp��+��7�ʝ��50V2�����K��:���˰�{���.6��� x��k��9�~��˗qS���D;��q�.uG?����1��p2\������w��~f8p��#���F̚�E�2/���x8�C��;������@CX��l�o��|��ë�_�z����p��5�G'?�8���Azo`��q7,v������C�����BjLGj�Ó�@�¥?>�Gh��n0��훻�������3~}9���D����[�i�{n7��og0\�H��{�m�b`VßW�s,L���@��0�_�n��@���ﾆi�g^'�������a �}j'��֞���|&����v�����b����1�l�6	���@چ�l���_�c{������� ��9�l�=;    IEND�B`�  Left� Top� Bitmap
      TPngImageListSessionImageList144HeightWidth	PngImages
BackgroundclWindowNameUnusedPngImage.Data
{   �PNG

   IHDR         o��   sRGB ���   	pHYs  �  ��o�d    IDATx�c���?5 �A��4jШA��A AGѡ�P�    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  RIDATxڽ�Oh�PǿY��m�?�X*�$�ju0�0��NE�e=젠 "�/<���@<x��AAA��@��)�2�Iݴ�Y�u��5͒�ϤiC_�i�U���x������X��|ǚ���4Vr��P`�P�';v� \{s���~��P`�1 ����aX��S#5t���#��Lр.����3#����b�^��Y��es�?���1	� �����	G���*H5sM��ү�!��p8yt����zT?A��ЧCE	Hf	R"�	D�`a�*�bQ`wt�>x�nv�yeL)�hQ H
z敊�]A|n�ضn����ي]�A˚1�S�^�����H���6;����v�yjuIԍ3+6-W��%,$�4`��-�u�>�:t� ��(dZ���\���/`ݰ	�g�ec�sY��F5��ҩ$hk��{�1L-r���5M>8!��Kz/>]�qI�{� �0sf��5��m�,� �e�ml�>S��7E)��w_S�_�D��������n>��i횓��"j�KmI��qXZ˛Q5W� ��{���h�����w�DM�M�|����/�?�f�7.�M([5'    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
<  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-�з Dlj��f`b�d*�ɯ���QTX�/�- ��̸_��CT\U*��o���������<
"��M��/4�\��U5��a������=/n� ���s�j��-�5Q��Ex<����Ӡ0�-���;�Sk�\Z�W��O�eT�x,��]������m���**���_g�m`���9A�=����
�@��Ud8û'O>��`�qm����?�f�;5r���`�;��2Hh�2H�1���T|��?n�<�����Z����a0�of`b~����+���/~�6�w/^�-P�o��ph�&����>���_��gd@/����2\�����_���X0ܻ���$ ����8��X�|~����ݗ��Ih��9e&6y]�??�p-�� �]����S|k�-��gP0�b�ef���-i�Gc�si�Y����G��=Y� �֑L���?�'ϒ�+��oóG�;z�����1���1��r�Fl|�b~�e8}����G�`m�V�/��Ϡe ��o!l���wNm\����q ؂�
���E8����H��'>0<���Ŀ�q/X��V�������"���?v��3������lj�}���(�@-����+�*��_� %)c�^c�    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
9  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-�𰀑��as�����@!T%��0�������)��`K�4�p���f�Jf(
�:���⩫��8�b	���������f	)8�[��aA���������+�0�X��K5���i�L�|+�P����&���b��v5T�4�#��sfaZ�]������8°�?n��s`Z�U������d�S~�ܥ�x.b��i�>��{߼՘x�Oe���V���2�w�F,�3��v
�&�|��ў��0-pϪ`���2\#���gٞ�{0-�e���:C��#Ďﾁ%�u0�����A�Y�}j7�֞F��|�k #W#�=��>�d�]�W����l�6	Ղ-��G�RVT@���T?��[@K@s 	�E�35�    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
o  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  !IDATx�cd�1`��
1�o�Q����n3*Į���D�Wm�� �@HT�&�{�b��rG���E����P+�M.�s?�,�6Ǐ&A���	b��Y�`�Go�� k5�|B �^/m3Ăs3|h���-NM�l=qL{[���0�f�[!��MX�B-8<�,���0�n���O����o�X��ϓ&>p,��`w�X`߹�`��H/���w-��`{�;M|�Y�b��N�/���Jx�� L�W9��p�lhb��#��Z[p�V��7i_��� �\�(_��    IEND�B`� 
BackgroundclWindowNameWorkspace closedPngImage.Data
{   �PNG

   IHDR         o��   sRGB ���   	pHYs  �  ��o�d    IDATx�c���?5 �A��4jШA��A AGѡ�P�    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  cIDATxڭ�mHqǿ���ܚ:��T�iM�퉴�
+
z���UaT�/*�=bM�QV�C�*����h>�����p�6==3������������{ ��(;v� &�G`�S�?�Y'(?~��(?�Hӻ�Q�v��/����P�K��@�Y�ڪ
_u���n�RE$�R�U�ʘ ���U��D1� +�q��|��������b<�x�9ԑ
�4105wb�f/������ ���5��=��+�8�� A F����s@�L������׍0�8H��3 ���r���B�v�1p�v��Mϰ!kʊs`��`1 #E""F�:t�=E��.�4�)Pn<��L	/6�5�Q�Cƍ�F�<��	�`"N*��=8]ۀ���xQwy
��"js56���;��w01�F���шs�;�
W��p��x�r{�sȆ+�aw��q�I�+��u��_�3mz���Ґ�2��1ĪáR��C� :>��氰�9������M�fG�䌮C	��,F�]�zM�
�m�$�r�X����'��T�k�t B���DE�A[V��DQ����萰���O��i	�05�^���ٚ�;&3����__	��&��D��X����C �aa����\�h���[��_�bltDP�G"c�-�	9 ;=�0�~���,]��� ���uw?��6!@�P"���܋���_|��xs/�v!@&�#�ЃE	O���.�4%H%R�[[�$��V0F Ir���_�#s6>�o`}i+��.X��'�E����p�?�![����u�?'q��r�v2gh��Y�����C�P ��5��@_��>��{���M��e_����X4G,ܢ��?m�]�Ʊ    IEND�B`� 
BackgroundclWindowNameOpen new session closedPngImage.Data
{   �PNG

   IHDR         o��   sRGB ���   	pHYs  �  ��o�d    IDATx�c���?5 �A��4jШA��A AGѡ�P�    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  �IDATx�cd�1`����^ǙYX-�i��?�O�>��j��eu=��<T1�#���7/1�>��n���6��9�T� <������)i0���CBKݻ�j���
úE�bAP\Ó�wP-��Qdظt2U,���ex��>��r�WL���Y/�?B�@DL�a��YT��+4��ͫg���3�X;�*x'3�{��~Aa��R�׀x���ߢZ��'��w��X������T��yl[N�"�}��já���b��{Ï�P-`cec�������e��������V}L�jUe���/�v�G��U����>�՚�
GI��?2�ލD�ũl���"����w����D������UԀ�߿�"�.
o�-�r�#*����D�(AD �D� i�b��:    IEND�B`�  LeftTop� Bitmap
      TPngImageListSessionImageList192Height Width 	PngImages
BackgroundclWindowNameUnusedPngImage.Data
v   �PNG

   IHDR           ��   	pHYs  �  ��o�d   (IDATx���1  0�_�P�A�h�Υ�@ �/��_���    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
n  �PNG

   IHDR           szz�   	pHYs  �  ��o�d   IDATx��kHSa��g�Ԗ�׼�d^�L������!�nE�AEQ}�>DQdBч"��.�Dbּ��f��es����t����ީs;������}w���y�K���`rTU�[�І(�Qs���N 9*kҺL�rT�������F�܁B���*���h���V4��P. 	�4H7�Gi��k��e`0O�c���:������z����S�%YR���A����j�4����׭&�%$C^x�)O=�[6f�ر��u8C�N�g���A��W"��*��$n�rg0�>j��Fz�q`�0�՝�.2@T���װ-E��y3�u��d0ƚ��;X��ߜ�ρ2@d�ZDn��<��i��:3k:2�Ls�;�N�W'��N�X��7�Q!v?�l샫Pk��څL5��8�~��"�Wr��"��Yml�j���.��Q�ώA;4H	��b�-l�9�5�V��`��-�خ��G1�ՐV��C��ҢD���؁���خ�Ǉ1:����{H����K�L�o��j���nl��*0��*.�����p-Vm`\?FX)D��*��:���^L�d�� 9�U
��n&'d ??�y"(@��R�LF2�L�[��hh|�y� �H1��n�c˕�����IĢe��Y�6�+YN�`�r���3��J�RZ����3���oI �Y�� ��|�����f�^�T67���zo�8E�S��GM�K�g�v� ��ZhQ�����<��G �� }��0?ϡ    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  oIDATx��YLQ��QY�P1*Z4JDq�Ke	�.DB>�+�AM41�d���B�7L4j4��1FISæDD@ B��UKC-Pʴ�-�8�s[����M&s�̽�|�9��p�σ�>�*B�r��2�NaO����P�ax|q��čN'��`Nn�����[�5Z�̘<�0/9j��Ju�."Z��<�D̓���?5zL����̬��\����1�XE��@%f�QAG�͇�hMT�)����
Pr�:4@�~UX��1�ؾ;b�~k`1�a�!�����3��axePb�ɲ��<)Nu�팢 6��Y9X�2�"������C��!���]��������<.�!'BMl�憹�Ct�1�IL��@��b��p���Y~�O������RQw3G�R 2<hi䐰�� uQ'WH����`}������|Hs��M����@��kd�'x�}���4�Ȼ�lfI[������:W��P jR���I�|�:\�rO��O��c
�"Y&���+�7�i���F,]����b��=��Zf�~��w��9P����$o\
@�a��t$��@��ʬ���"K9����nE���F��Đ�S��!6^	�`	�0t���7=�h�����Wd �Hkw�bJ?Y�`�a�g��I�����Y�35��2�	�)����s�k����7�����p��cЭ�Ud�L���U�� vIT@�NbS_E����K��.nT��3�����K,X�
�6f�N@z�?��ͣ\��)9�L���qPΌ���%JA�LpTVm���s���f�y��|�	�^���s�R�ǿ˚[o0��ړ��3?��/�����w�Ǭ�E�v��� ? +L~?�
�    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?�@�Q�: � FFF��",r{�α¡�ȏ?���~�k6����E�[�>�D�*���G'0�8��ͯ�q5���Y֜���ih*#+'VͿ|c8�z�߿_���6<;GUln�����#���׀���0\ݷ�� 8�[�����;'�k0Q`��@0�t�}�Mpp�%����P����ghj��v��.�����&$��Te�3��J�3|}��h�It��9s�;��x=���;H���Ca�܅��Y������8!5D0���]B��~|ޏ�@�����+�;�#:ï/�������yk	8 �����$?���H�9�����Jpc���y��;�=���Ϗ�DY���ՠ����E�yަ��q9`~��'3����aB����=�~��:��v�ϧĉ�}�@I�[�����&V�����`�	t�oTI*Y�v? Pfi�R��l�6	��>�<4@{���<��ꀁ�  Iӯ�v �	    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  �IDATx�cd`�8� C!f�- O�N��|�8P����gE����i��0 ��� s�8�Ε����'D|���f�;����bH���H�8.����������%
�7bw��y~tq�F�&��6‵Gn�h�Q'I���J��+��:�8pi�/����-�j$��0�zi��;��L_���A:���fo:~E���*I� L�Q��83͇.!`�����z��[O����B�$q\ ��,{+v���M�����c������h�4S!I����݆�G&z�%l�q8���v�A����
I� L�]����K8n��}}�9{E���2I� L�S���K������(�4�ۗ����]�tq�g�N���Ix�cs�@wL
�:  ��	0�,�    IEND�B`� 
BackgroundclWindowNameWorkspace closedPngImage.Data
v   �PNG

   IHDR           ��   	pHYs  �  ��o�d   (IDATx���1  0�_�P�A�h�Υ�@ �/��_���    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  �IDATxڽ�{L[uǿ������UE��enlL̖0�f�t�2�fF�4Ӹh��i`1�f\�9ԍ9���]��?�1���
�&���װ`ˣ�R���߽��;�깹���~�����s򻗂m���]b?�i��)���Ǆ|(_�y�^}H��죦N5�={�({�d�ÙIƣ+ĵ����;�M'�t�JuTJ'�$_:���P������[) y����<+̄�0��7O�j��<$�(��J�'Ln�u�ʝ��y"o��Dd�(@Qs!��8�*��ՎР@���f$F�b�d��6i������r&9-T�k����<ˁ��E :`�e�;a��iD�KĜ�*��4|��5�Uu� �R� )z�uR.�v���\W�O؜�-E�0Yf�C�J.��fFF�������M�1N����Y�[ؙ/q���%�	���WP�x>cø�ĩy���Լ공�� /�Ey�d.0���v�����s�N�Uؑel8�H�Y������ߠn�Qs���u@\B
�K���,1_hQ���Q�Y�ʊ"�n)h�F�T����[mv8N8���u@��W��Q(������7�`��]�u5�YR�!�� ET��2��?�˭�\Y�?8��7l�D�&"��6����^M���H��iz�0�k��d0XH����%��Cp�W4:h��0���p?4�-{ 2Z���'Q��c���19�����An�6�t508g��sh��8�-Z��*0�r��!a���X��� kD��#٭�؝����Y�P�&E�Ά�������aa���((w}��D�&c��d��i�{��	���[0��%�J!�G���3���F e�'Ȋ�k>9�`t���҄=���Ds'������� �k��R#)��FL����^؏�	�0��5Ȯ<�9ť�u����<�$�L� ��A�{�q�E=���	L�M� ��r�}��O~�l/,�0@@�U�>�ԫ`��H���X��� m��`��
H����_�u���aw���d����O����I�ګ-~|��m�����cܧ�+sN۪��X�%��
}��%��
 #�A�[��W�4�����s�m��b����r���+3xs��o	�
���}Y �Kw,�&h?~yE �`	�����j�I���    IEND�B`� 
BackgroundclWindowNameOpen new session closedPngImage.Data
v   �PNG

   IHDR           ��   	pHYs  �  ��o�d   (IDATx���1  0�_�P�A�h�Υ�@ �/��_���    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  7IDATx�cd`�8� ���{	�Mk��g����陃��P`b��WUS����}��3��2�����%5]���ijyDj%ý[�N�ʈ� -�Us�hꀰ�2�w�aw���Ú�=4u@Hb	ã{7�;@VA�a��>�: 8����[� -�°~��: 0����;� )�Ȱq�d�:�?:������ .%ϰy�T�:�72��峇� &!ðe��:�'<��Ջ'� "&Űm�,�:�+4��ͫg� $"ΰc�\�:�#8��ݛ�� ($ʰs�|�:�=0�������/ ̰{�B�:��?��ㇷ���'��w��:��7�������ǰ�2�:��;���O�����p`�
�:��3��۷/�����ph�j�:��=��Ǐ������`kcMS>r��ׯ�����JKY�n����~���� P�����.M�?�a6�L�1�g�fdd��#��҅�Fi�H
j����?�u�d��r���%Vܸp�� &�+@JY���_Xղ���]&6J�_VQE���X�bSK�9��ɏ�2��ؾMTq F� (�Z �5�!���y    IEND�B`�  Left�Top� Bitmap
      TPngImageListActionImageList144HeightWidth	PngImages
BackgroundclWindowNameLoginPngImage.Data
E  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?-#��V!_Ffƙ���0�������|T�~#���"��R��Tq��?�����A�[i�����E�
J�|�C���6����[��a�Z�?=���~�[F�R�"p�G<o00!�A��f�����T$u��
����V[Ԉ6]��+oQ-��+>�wL[lR%�t=/��C�@LC��d�0m�AL7��1t]�c���N������QU��S�w���Ze8�ŷg5��.�=��t=�o@� �Lq��t�=x$ν6�a�R65����40��Z ���p6�>Q�}��y����Ͼ>�����T���B�@P���\��#��/g���_���-W ��~F�@@���|�C�- Fx��Z�0��K����_P-���f���� zs���P��/� ��5X$�?>��j�N/%<�G�̋�x�����[ �?���j�'n'=ax��)C��l����T��d���W�Q-��+���L�̖ӝ����V2|��;�������\����j�30�=S��HG����OT8�����g>ӚӉ�������vV���dךS ����6.��f�^�P�h�,���R�ڽ�`��o��Lf6&)&&�]��������*��>- �2��V��t    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   IDATxڝ�kHSa���9o�CWy�:sMsy)E�@��Aj6� D��}
"�Pt�ԧ����@"�6CĜ������릸�2�b��6��u�����9��\~�{��	д���!���o1�'�&ǧd�a�_3鏱�0/T!7���V��7��H�q�	ʗbf���78)Z8�w½�
�>YX\�,��|]�p�Yf QQ5��ᢩ���}xbR����[&�� �7<i�<�g�)�A��x� ��ð�-d.1�N�[�(ϣ8��IeyA�=���,���� �����ߦ�Y.=�䮿P�{�HT�aGOPUm͐ϥaܫ�a]wY�΀�;�lv� 9��+�Z��+F|�,�,�F�am����H��J�n�ODi9,�_�u~fDi��8�u���+o�@8Rhl��e�̇�n��{��Y�XvM�A���.�&)4�ЄD�u��ej,��7X`���֣�e
U.�ܔZ��;)���Wy	��bl���-�բU�V��9Ϧ��[�jتP��lx(J)$�K��|×f	�5"����v>���T�Ŷ�)&�W��B�89�13܇����䠺^N�S���Z$�gQM$f�$���﷐�F�d�}�B5�G�rtT\�y���/�!��	-	�����^[@�t
�
0ji��g��X%<(�2ė�ÕM�`"���rĳ*��2�3Pr�Z�E�� 	��m?�s7��{Ӟb��E�� !!�trm��g�ѴfQh��� -���@���:��P�fSh�͸�����<~�]��
�k �nw�*�y�    IEND�B`� 
BackgroundclWindowNameRenamePngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  =IDATxڭ�kHSqƟm^��YW��e��T����vӖfe)*)����0-�BҰ,�S��%��$#����ּΩ9�l�L�e��#'�yk>���{�����?�A����	d�t�b��_�1�pǖ�hg�=�D�Z��;M���gc��c[�v�m����k�ԧ*�$B�t��+��=��˻�kS�R=�5H����]��\y,4���f]��V��q�_,AT��H`��֥��z�J��ɕ���Л�Sz���3(��o�d��Ԑ���A:R�q�0Яr-{x��,@�D��w淸nc[?���CO;��
���������t��;����ցaTcXل���7�\dz�q� e�N;�l[�R�&�s#�:�eZ|�~�4E��s��n]���7��Śm�^	��-��i�ũ�G��3' �փ>ًV���B�\�)���ZuP��m��^���gے�}�;��RԼV$�n}��Y�`����y�#�ڛ��0��W����N�d�gu�\@Vn\&w?4M�nk��jo(+�ݥ E��S���.܋�A�a���1m��9PhD� Λ�<<�`p�R$".�s�5��A�i)�_���1�<�b�C2�ڿC$.��?-��� w%T#ZrtM���S�uK!r�ķ)t�
X.;'��s#�(@~�)��~tM��� �%8��h�p9pkF �G�ROR�3��kZW"q$��L�x��M��lN�Q���I��A�?�
�ǐ~�y�pp���1-ҏ\O
G|V�V/G�W9�3�)q�IHw��9��"=)@V�9/�FI���G3G? �X$�@��    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  OIDATxڵ�mL[e�������A[
�!.���-1�,ƨY41j̒}��׸����Ęh��l
,d1�,fY�,N7MP� Xpcl��F"}�Ͻmoｽ>�[i��a�[O������Lӄ�ih��8?�_P6*v��Ǥ�Η�:i���s =��i�^��z�� ��D�[�m�@tX����c��9 K�a��w��@cc�'��_�_]O�K��)�tK[����`p`DSS��S��2�nAx��`�ڽˇDQ C7�`�Q�v@��[K|�P��;�3.W`,�/���gz$ib����2ɩ��CW@��/���)�$����G[��(�O$�p�TU�i:�D]���e�3�m5|q�+#�H�p98j��sE9�)�$�+r�[��u�t�AUS�?|���щ�M>.:��mSM�����@����q-�������o�#����[�e�4.�����~�?\��;E���E�S}�oE�7���ݘL�F��-	����E�a04>	��r8���K��T[���RMyYEUYIƿ��az~�*� �!0�&oN�|�$'?��Gk�纈��\Y⭭�\b�Ά+��L8zv�O�{/���@!'���]m�Y�3s0���G�x*����Tt_��]YU���o*����,�9�0�j6��bm�g�Rv�r��a���u��� �1�W�s�^��L�2�Y�?b24����|�	�OY�8�_]���.������y�Ñ	�'���P$d"�H3�f�4����(�%����goov�3Ax���S>W!S�2�p*#�EE׍ݝ���.�?�٨�}�B�����Ht�ԉ �;�z$a?�l'wHHX��e1]�_c�n�Cd���cފ��I"%�At�1������y �x缿��ur�HCPQ�OX�}u��4��4��&�h�Z��~(��ë R;��B#���I+8�4UH��)_�F��ʆ�k y^�����d��3��z`}�,HM�7IiH��)Ga��F��~��)Ct�izH�4_ ��Ι"����Kv��뉯ا���B̏`"����r}ݗ�Q##�(p�@�oN���iL�eX�    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  -IDATxڵ�yHTQƿ7N�W��ᒤdY�(�ZZ
j�hR"������FMA�F�e�����V*ZF3�K�KJ�D�V�:��8��̈́cΛt��<���~�=�>���0�����mB=!'����Sؙ�}5`�ǁ���!��k��D�?pY�)��YGb�T����=G�9�M���i�Srv�]�fL��/�[v"vF�
d�`3��m��Y+�š:@9����M*�K��(I�(�*$���� ;��eA�Hm�|�5�r4-Lg���BS�'d�⿻���T�r���5�k��;{�� ��j�(��_���5��s����!*�#�Ƅ��0e#��]E�E�q/���3.ʹ����D7�sT���h\\l4��hn1*U�{�������� d˞h�����W+��l|8�-1VB�\I�K���Bd
ȐH��o_a�8m��6#pc0V�;�P�����6GsgZ:���5�G$h��]0ֽ�X�T�'{�h���6���zO7>���0��;�H�jJ%�4������j�9q ːz��A�q���ǂ����ǻ������B<p��D�k�O�B��s�j/B|��7r����'��L)����X� x�VX�!��l%�so2[�`T��(��K6� �6�X �������sO�W�ʂ|�Π 5��h���2��砐4L��#�����?���qx&0~>�	������@����W�N�(�<�j��A�	�Uf�3>!�P+œ
R�B��^�<�Iƻ&�C*�e2 ��/�Y#u��{�t���~��Z����    IEND�B`�  LeftTop� Bitmap
      TPngImageListActionImageList192Height Width 	PngImages
BackgroundclWindowNameLoginPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  (IDATx�c���?�@�A� �F!9Vv����m��l�������G~�������#(����u��d`dd���@�>��������*�9�8@�C觴�(�,Gv���ݯxǎ� ���"4��^x�p��-#����;�L���O.����������d�R{v	�$u��r��&Y�#;�z�:����[����j�q��`�r�*ɖc����;���j�	�;`�b�
�������� ���'!�����a>���BÇ��	: ]/������X9|L��U��?�z��~��a��x��^����"*�D��{p6���q�L��%�؛;�;@X�8�	���� ��3�������d�o��p��\�و�D9��z�
%4`��P���{�	��x��E= ��� Zr��G�Q�1Z� W���g���+:��l����; f��Ry���_�;�_���B�#�-Y�|�%
`�,���}|���$����b<��@6�`��p;N�����x%��r����p����������Z��p��/�aw �1�\Nz�u���� _7-g��`^Ǣ��/�F	Vp�p`5�J�S0�3GL���fh<R��;���������\B�p5b��,iR6����p � ;VC��?�Z3�Hv 6������ ~��k��(n�hMG8���_��΋��]a�1d7�V]]�P�.��3�q���KR�����9@�'+0h�,���o0�堎	3+�#M��������0;&�5(0�  �C�zl/�    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  YIDATxڵ�{LSWǿ�R�RI�aiy���,��
cLQ���۲�%Y�����,[�ÄefK��dd.�13*���q�:�YH@�R�B�j���g�Z)-��u��=�����9�����R��^-�s��G�6tR�T�i.��1�R��8s#�k !�n�/w��ڵt��?WO~��Jv "��kd�]d1���k�C�@�;�3�h��	;�TQ��Zq������`tk�o����Ҍ�HN�my��ҝ���3��'	?y�sLO����㭺X�0`Vc��g�Q	��z6h�xK-��Iv ��d�7���H��l�@��	n�w���)f��� k���;���&l��y�{0=�@�nT��A�6��0�g��'���ld�Vl�8n\�Ϟ�ߒN�9 �N��9@I�.������KDގ}�pc0�����(���j��S��b6E���(gƲF�_��m����4}-��]1D���]ݰ٬��|�V΍�6o,�)H�y�;n�kq�\#~�ѿ����V0���\������qyq�eo��֧���o]ù+S�McF�C��j�`�&J6s �y <����t��}�g��j��N��r|N���7J��jے��Z����t�q���X�(�w�;SNE��-�{-LI�tG{������jq���4-�숦�(8$g*�'�ąG]mPj����H��ˠ(?�pT�?z��^l((���a���K�;��{�DJf���jF��(�Q�����b�a�_�eN��1�u}��k@(F��jY��(Kh����	�hI�w�d��I���P�X�j�@K/<g%�G���O����2�E�7ԏ�7q�/.�Gt�Q�Um�L�����{,�|e8���C�b1�b_
�&�~��Gզ����b���%XK׋�ؔ���Om���:F�X��˖����
���v�s5�UTc�Q�N:���+��5���q�7�4r�SbF��@�h�y}Uc�㽄��oʤ�!���$��}|Uc��DŖ� ��ܪ���gAD ���Z��7!�HTt���뵏}|�T�E��7��R��%A�e�?4�B-I~�3    IEND�B`� 
BackgroundclWindowNameRenamePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  RIDATx�ݔ{L�W�_)-P� �r)�v�6F�$�faSaen�A�Dv���$e��"ddW�.�	�1↗m�f��eQ� �\W
�@�7�Th��>C�mR�������=�}����x�!�������`�������% ��������#SӐ���'�SY{��%(c���^E���I���n��1��,�nء�)�aRIK���t�;����Õ�rZ�d�xyW��q�1W�8�?~n�h�+��6m{S�����E��9Y�~�tJr��2/6~o��H٧�q����ӞE8Kzz���w19�^,�~���c�jT�s�3r$����C��*c_��`��/���?�ޯ}Ϙۻ����.����-�@}w}���Sh�*0�o�|O�L�/�ĩw6Y��&PE���}Ek܎�N
f��4SJ�D�Vr���/X���{tM�ڃ^��C���Z4]?���+z��	ԑA၏�K"�#igLF������d�� f�08L�$A�r�5ŧ?�t]nd�^&F�m#z;����^�˜y|{��/jC��~ �?T7�Q����
��g�uμΐ�\� ��5��]�˭�`�N-�~��ЩB�I�ڡ�����]<#A��@#=	y���۷��N�3�n˃�ZXlTm��A��6aRu��� ;��'{��y3)�}m��ba���j���g�`6Mc��C�j5�V��q��]�S�{�5�~oZ.� $L	w�z�h�۾���4���n<]Tn+Puh72>�@T�m=�~���j��T &�Wn1�#�,E�����:��7�,��7f�����ٹu���1��
�S`�/A�g�ʄ
�-[i���|Eއf����ٹq�A~���C7:��*�'�{�n8ű8��1�x��
TMe�h��|	���ń^�Z�^�'Ƽ����v�4�� US��"���O�02���ͅw�F4����F��}��'@�Tʊrq��%d&�!q{X\��T���ܝ3��ՠj*v��A��b�"�86%��Dαj����"���M��$i����(pk�,������`I��������G�?�e�0�J�Q    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
}  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�ŗ[LSw���sN/��@�e3N]A�RD�K��%��OK�3�x�q��Ӳa����MA�|X�qƩ�,�ѭ���TJ��\ZzN{�o�]�����������~������
�S� �a���f ����vI��O���ʲ�#G �{@��i��K�$~C�Ūih⥳Yb�58�VVn�{�}�>h���Oj�;�������Zb�7W�ʊ"7���4��q�f�U���\�ܡ�d�a'ϟ^��C��W�_+*��e˖��������v�yz���6���6��LL<��گ˲ys� �>_�-4�:N৫�J�E�����B{�Mx0�����ߟ	��M�T��Z�i��y}�����(6풤���f���OتJɂ���Ed���y�F�;��jx�Q��%ߔ��Va��6E�����Uu�Apf}s�ݮ#����,/�K�w�xr�x
Ͽ�@H��-��8��Vn-I�m>xo�{���h�f�G1��A�����X�J���qC�{�)�N;$C4h,�R�[�f5��4�����C���<?����n�O�s���=�DT�nQ�$�[Z�Sʠ;��d%0�!�90�{�.%����,,�G��!h-I$�F�v�o�J�6�c����c�jq��Z�KXM�$@:7�[G���H�g����+fĎgb����Qu}��� ��Hb���U��<�I���7��+�A��$o�x�= �����|Б)X�0�	�-�S�ˋu攨��I��_��q�%�Ueˮ�t�ȼ��B��meK�K�r�>'�B�軫N)�w��$<F���R��?^^Thz!Q\R$��10�)��.�0�,��*Q�]�Z
L����{$�~� �&��`���^ıY��ahQ��Hc�(�x& -,�6�᧪�
ɂY�I705�#�r"���t� ZYz+�i��-*č��bL�kl�V� OI�	�W=^e�a+G��b��5�|�����-Ԧ�ҥX!2���H�x �o�G�u.D-�9��Ԙ�@�l]�����d).b�#r{-�2�>��5��Fd�fg(��9֌8�'�Ts@��-���]n�݌(\�߆2$U�B� �݌��H��U�즾IB���:E1k;na��z~p-�C��/I���N�^��HF��@�G[*P��r��-1�!\����,� �iQ�V24��r|����
gHb#Y�^�k&��ܫ(p3�\8���e�IPO�S2?�;��d�qT�#.��ttA�>�D�3��
��Pzi.�IO��k8�9�F��͏ b���:�FN����� ��5�!�"!�)�#Ve��x��|�'=a0�h⼕$L�����%����D& V�8�RU�ԭ;�O5�����ί���Fd�K������eH@�F�fǞ٧A\D��" ���n��Ҍ>Nsi:g�(>��Ox^�/��1��k�    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  "IDATx�Ŕ}L[UƟ[��6 �D)Ω�q��d�L�bՍJ�)�,�0�|S���0����u��tȇ�E��f��+u3c3�0C�
C�A)Ю��^ﭢ�v��+Ž7M�9������y{	���AudU�$Tyf�j�p��b)2wU�4S�G��� ��2�	�}��4ay���|Ua8��e�i4:1)�����?z� ��z�v����DF��QX��Y
��H�,_�nr�)��Z2 ��ɵkבJ��դ��� :"C�6�t��UѰM9��C��僉!�(�*Vm|�m[�HR���x1�݈����"��D��Y�yi��F���@��a���%�%�ۯ�Y�Y:���PV�����r΂�&���[_F��;0����U�6ǧy#@�x��)���`��*-핸r�ဪt���� �8��<_�N���90�����uي��0��k_�8V�(	?�^�!��X�=���h���u:�T�7�۞�wUt����qw!�����8���݉�ӿ��ٞ}_뵻���\���r����k8��Ͼ��c:��n�+�ぽx%-��[�$!� ���x缘�׿5u���_{@���b�MHR�
dmUCB����I_�{WF!r���1��ka��K���Ǉ� R����p,�+)a�<z���P=���~������ѵ���� �����&��B`�����{��[�ԧŗ?��3�^�K�H+�\k|l� �x<n~φ�Ժ0��&8&���Z��6#���(��9y( @��q�I� n������`K�w�n?q{�R�1�6p���
.{Kж�;r���ڣ ޮ�k��!���h�5pl~��3?��~��0�5 (8���-�6[����X ��2x�]A���SuFn�My%�s���o��T}K ����ZBb7;@7��ٯ�t[��ki�?��t����a�W���ϵZ|	��"]�-�wϏ�Tp$oR� ��D��3����K�f�MS��4��h<\� ���˱�A�I�=���N���ʂ�.�    IEND�B`�  Left�Top� Bitmap
          TPF0TMessageFormMessageFormLeft�Top� BorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionInformationXClientHeight)ClientWidthFColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterPixelsPerInch`
TextHeight    TPF0TNonVisualDataModuleNonVisualDataModuleOldCreateOrderHeight�Widthp TTBXPopupMenuRemoteFilePopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�TopP TTBXItem	TBXItem23ActionCurrentAddEditLinkContextAction  TTBXItemRemoteOpenMenuItemActionCurrentOpenAction  TTBXSubmenuItemRemoteEditMenuItemActionCurrentEditFocusedActionDropdownCombo	OnPopupFocusedEditMenuItemPopup  TTBXSubmenuItemRemoteCopyMenuItemActionRemoteCopyFocusedActionDropdownCombo	 TTBXItem	TBXItem72ActionRemoteCopyFocusedNonQueueAction  TTBXItem	TBXItem69ActionRemoteCopyFocusedQueueAction  TTBXSeparatorItemTBXSeparatorItem9  TTBXItemMoveto1ActionRemoteMoveFocusedAction   TTBXItem
Duplicate3ActionRemoteCopyToFocusedAction  TTBXItemMoveto6ActionRemoteMoveToFocusedAction  TTBXItemDelete1ActionCurrentDeleteFocusedAction  TTBXItemRename1ActionCurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem82Action#CurrentCopyToClipboardFocusedAction  TTBXSeparatorItemN45  TTBXSubmenuItem!RemoteFilePopupCustomCommandsMenuActionCustomCommandsFileAction TTBXItem    TTBXSubmenuItem
FileNames3Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItemInserttoCommandLine2ActionFileListToCommandLineAction  TTBXItemCopytoClipboard3ActionFileListToClipboardAction  TTBXItemCopytoClipboardIncludePaths3ActionFullFileListToClipboardAction  TTBXItemCopyURLtoClipboard3ActionFileGenerateUrlAction2   TTBXSeparatorItemN1  TTBXItemProperties1ActionCurrentPropertiesFocusedAction   TActionListExplorerActionsImagesGlyphsModule.ExplorerImages	OnExecuteExplorerActionsExecuteOnUpdateExplorerActionsUpdateLeft�Top TActionRemoteCopyQueueActionTagCategoryRemote Selected OperationCaptionLadda ner i &bakgrunden...HelpKeywordtask_downloadHintB   Ladda ner valda fjärrfiler till den lokala katalogen i bakgrunden
ImageIndexk  TActionRemoteCopyFocusedQueueActionTagCategoryRemote Focused OperationCaptionLadda ner i &bakgrunden...HelpKeywordtask_downloadHintB   Ladda ner valda fjärrfiler till den lokala katalogen i bakgrunden
ImageIndexk  TActionLocalCopyQueueActionTag	CategoryLocal Selected OperationCaption   Överför i &bakgrunden...HelpKeywordtask_uploadHint>   Överför valda lokala filer till fjärrkatalogen i bakgrunden
ImageIndexl  TActionLocalCopyFocusedQueueActionTagCategoryLocal Focused OperationCaption   Överför i &bakgrunden...HelpKeywordtask_uploadHint>   Överför valda lokala filer till fjärrkatalogen i bakgrunden
ImageIndexl  TActionRemoteCopyNonQueueActionTagCategoryRemote Selected OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionRemoteCopyFocusedNonQueueActionTagCategoryRemote Focused OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionLocalCopyNonQueueActionTag	CategoryLocal Selected OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionLocalCopyFocusedNonQueueActionTagCategoryLocal Focused OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionLocalCopyFocusedActionTagCategoryLocal Focused OperationCaption   &Överför...HelpKeywordtask_uploadHint3   Överför|Överför lokala filer till fjärrkatalog
ImageIndexX  TActionRemoteCopyFocusedActionTagCategoryRemote Focused OperationCaption&Ladda ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionRemoteMoveFocusedActionTagCategoryRemote Focused OperationCaptionLadda ner och &ta bort...HelpKeywordtask_downloadHint\   Ladda ner och ta bort|Ladda ner fjärrfiler till den lokala katalogen och ta bort originalet
ImageIndexa  TActionRemoteCopyActionTagCategoryRemote Selected OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionBestFitColumnActionTagCategoryColumnsCaption   &Bästa passningHint6   Bästa passning|Anpassa kolumnbredden till innehållet  TActionGoToTreeActionTagCategoryViewCaption   Gå till trädHelpKeywordui_file_panel#directory_treeHint   Gå till träd
ImageIndexLShortCutT�    TActionLocalTreeActionTagCategoryViewCaption   &TrädHelpKeywordui_file_panel#directory_treeHint   Dölj/visa katalogträd
ImageIndexLShortCutT�    TActionRemoteTreeActionTagCategoryViewCaption   &TrädHelpKeywordui_file_panel#directory_treeHint   Dölj/visa katalogträd
ImageIndexLShortCutT�    TActionQueueItemQueryActionTagCategoryQueueCaption   Vi&sa frågaHelpKeywordui_queue#manageHint'   Visa avvaktande fråga på vald köpost
ImageIndexC  TActionQueueItemErrorActionTagCategoryQueueCaption	Vi&sa felHelpKeywordui_queue#manageHint.   Visa avvaktande felmeddelande på vald köpost
ImageIndexD  TActionQueueItemPromptActionTagCategoryQueueCaptionVi&sa promptHelpKeywordui_queue#manageHint'   Visa avvaktande prompt på vald köpost
ImageIndexE  TActionGoToCommandLineActionTagCategoryViewCaption   Gå till komma&ndoradHelpKeywordui_commander#command_lineHint   Gå till kommandoradShortCutN`  TActionQueueItemDeleteActionTagCategoryQueueCaption&AvbrytHelpKeywordui_queue#manageHint   Ta bort vald köpost
ImageIndexG  TActionQueueItemExecuteActionTagCategoryQueueCaption
   &Utför nuHelpKeywordui_queue#manageHintC   Utför vald köpost omedelbart genom att ge den en extra anslutning
ImageIndexF  TActionSelectOneActionTagCategory	SelectionCaption&Markera/avmarkeraHelpKeywordui_file_panel#selecting_filesHint"Markera|Markera/avmarkera vald fil  TActionCurrentRenameActionTagCategorySelected OperationCaption	&Byt namnHelpKeywordtask_renameHint   Byt namn|Byt namn på vald fil
ImageIndex  TActionLocalSortAscendingActionTag	CategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintT   Stigande/fallande|Växla mellan stigande och fallande sortering i den lokala panelen
ImageIndex%  TActionCurrentEditActionTagCategorySelected OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera markerad fil
ImageIndex9  TActionHideColumnActionTagCategoryColumnsCaption   &Dölj kolumnHelpKeywordui_file_panel#selecting_columnsHint   Dölj kolumn|Dölj vald kolumn  TActionLocalBackActionTag	CategoryLocal DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionCurrentCycleStyleActionTagCategoryStyleCaptionVisaHelpKeywordui_file_panel#view_styleHint9   Visa|Växla mellan att visa olika stilar för katalogvyer
ImageIndex  TActionCurrentIconActionTagCategoryStyleCaptionSt&ora ikonerHelpKeywordui_file_panel#view_styleHintStora ikoner|Visa stora ikoner
ImageIndex  TActionCurrentSmallIconActionTagCategoryStyleCaption   &Små ikonerHelpKeywordui_file_panel#view_styleHint   Små ikoner|Visa små ikoner
ImageIndex	  TActionCurrentListActionTagCategoryStyleCaptionLis&taHelpKeywordui_file_panel#view_styleHintLista|Visa lista
ImageIndex
  TActionCurrentReportActionTagCategoryStyleCaption&Detaljerad listaHelpKeywordui_file_panel#view_styleHint&Detaljerad lista|Visa detaljerad lista
ImageIndex  TActionRemoteMoveToActionTagCategoryRemote Selected OperationCaption&Flytta till...HelpKeywordtask_move_duplicate#moveHint0   Flytta|Flytta markerade filer till fjärrkatalog
ImageIndexd  TActionCurrentDeleteFocusedActionTagCategoryFocused OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesFocusedActionTagCategoryFocused OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionCurrentCreateDirActionTagCategorySelected OperationCaptionS&kapa katalog...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionCurrentDeleteActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesActionTagCategorySelected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionRemoteBackActionTagCategoryRemote DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionRemoteForwardActionTagCategoryRemote DirectoryCaption   &FramåtHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionCommandLinePanelActionTagCategoryViewCaptionKomma&ndoradHelpKeywordui_commander#command_lineHint   Dölj/visa kommandoradShortCutN`  TActionRemoteParentDirActionTagCategoryRemote DirectoryCaption   &Överliggande katalogHelpKeywordtask_navigate#special_commandsHint"   Huvudkatalog|Gå till huvudkatalog
ImageIndex  TActionRemoteRootDirActionTagCategoryRemote DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHint   Rotkatalog|Gå till rotkatalog
ImageIndexShortCut�@  TActionRemoteHomeDirActionTagCategoryRemote DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHint   Hemkatalog|Gå till hemkatalog
ImageIndex  TActionRemoteRefreshActionTagCategoryRemote DirectoryCaption
&UppdateraHint$   Uppdatera|Uppdatera kataloginnehåll
ImageIndex  TActionAboutActionTagCategoryHelpCaption&Om...HelpKeywordui_aboutHintOm|Visa programinformation
ImageIndexA  TActionStatusBarActionTagCategoryViewCaption   &StatusfältHint   Visa/dölj statusfältet  TActionSessionsTabsActionTagCategoryViewCaptionSessionsflikarHint   Dölj/visa sessionsflikar  TActionExplorerAddressBandActionTagCategoryViewCaption&AdressHelpKeywordui_toolbarsHint   Visa/dölj adressfältet  TActionExplorerMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHint   Visa/dölj meny  TActionExplorerToolbarBandActionTagCategoryViewCaption&StandardknapparHelpKeywordui_toolbarsHint"   Visa/dölj standardverktygsfältet  TActionRemoteOpenDirActionTagCategoryRemote DirectoryCaption   &Öppna katalog/bokmärkeHelpKeywordtask_navigate#manualHintC   Öppna katalog/bokmärke|Öppna vald katalog eller sparat bokmärke
ImageIndex  TActionSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint Markera|Markera filer efter mask
ImageIndex  TActionUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint$Avmarkera|Avmarkera filer efter mask
ImageIndex  TActionSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla
ImageIndex  TActionInvertSelectionActionTagCategory	SelectionCaption&Invertera markeringHelpKeywordui_file_panel#selecting_filesHintInvertera markering
ImageIndex  TActionExplorerSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för markering  TActionClearSelectionActionTagCategory	SelectionCaption&Rensa markeringHelpKeywordui_file_panel#selecting_filesHintRensa markering
ImageIndex  TActionExplorerSessionBandActionTagCategoryViewCaptionSessio&nsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sessioner  TActionExplorerPreferencesBandActionTagCategoryViewCaption   InställningsknapparHelpKeywordui_toolbarsHint.   Visa/dölj verktygsfältet för inställningar  TActionExplorerSortBandActionTagCategoryViewCaptionSo&rteringsknapparHelpKeywordui_toolbarsHint)   Visa/dölj verktygsfältet för sortering  TActionExplorerUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint+   Dölj/visa verktygsfält för uppdateringar  TActionExplorerTransferBandActionTagCategoryViewCaption   &Överför inställningarHelpKeywordui_toolbarsHint9   Dölj/visa verktygsfält för överföringsinställningar  TAction ExplorerCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionNewSessionActionTagCategorySessionCaption&Ny session...HelpKeyword.task_connections#opening_additional_connectionHintW   Ny session|Öppna ny session (Håll nere SHIFT för att öppna den i ett nytt fönster)
ImageIndexSecondaryShortCuts.StringsCtrl+Shift+N ShortCutN@  TActionSiteManagerActionTagCategorySessionCaption&Hantera webbplats...HelpKeywordui_loginHints   Hantera webbplats|Öppnar hantera webbplats (håll ner Shift för att öppna hantera webbplats i ett nytt fönster)  TActionCloseSessionAction2TagCategorySessionCaption   &Stäng sessionHelpKeywordtask_connections#closingHint0   Avsluta den aktuella sessionen och stäng fliken
ImageIndexSecondaryShortCuts.StringsCtrl+W ShortCutD`  TActionDisconnectSessionActionTagCategorySessionCaption   &Koppla ifrån sessionHelpKeywordtask_connections#closingHint=   Koppla ifrån den aktuella sessionen, men håll fliken öppen  TActionReconnectSessionActionTagCategorySessionCaption   Å&teranslut sessionHelpKeywordtask_connectionsHint0   Återanslut den aktuella frånkopplade sessionen  TActionSavedSessionsAction2TagCategorySessionCaptionWebb&platserHelpKeyword.task_connections#opening_additional_connectionHint   Öppna webbplats
ImageIndex  TActionWorkspacesActionTagCategorySessionCaption&ArbetsytorHelpKeyword	workspaceHint   Öppna arbetsyta
ImageIndexe  TActionPreferencesActionTagCategoryViewCaption   &Inställningar...HelpKeywordui_preferencesHint2   Inställningar|Visa/ändra användarinställningar
ImageIndexShortCutP�    TActionRemoteChangePathActionTagCategoryRemote DirectoryCaption&Byt katalogHelpKeywordtask_navigateHint1   Tillåter att annan katalog välj i fjärrpanelen
ImageIndexShortCutq�    TActionLocalForwardActionTag	CategoryLocal DirectoryCaption   &FramåtHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionLocalParentDirActionTagCategoryLocal DirectoryCaption&HuvudkatalogHelpKeywordtask_navigate#special_commandsHint"   Huvudkatalog|Gå till huvudkatalog
ImageIndex  TActionLocalRootDirActionTagCategoryLocal DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHint    Rotkatalog|Gå till rotkatalogen
ImageIndexShortCut�@  TActionLocalHomeDirActionTag	CategoryLocal DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHint    Hemkatalog|Gå till hemkatalogen
ImageIndex  TActionLocalRefreshActionTag	CategoryLocal DirectoryCaption
&UppdateraHint$   Uppdatera|Uppdatera kataloginnehåll
ImageIndex  TActionLocalOpenDirActionTag	CategoryLocal DirectoryCaption   &Öppna katalog/bokmärke...HelpKeywordtask_navigate#manualHintC   Öppna katalog/bokmärke|Öppna vald katalog eller sparat bokmärke
ImageIndex  TActionLocalChangePathActionTagCategoryLocal DirectoryCaption
&Byt enhetHelpKeywordtask_navigateHint1   Tillåter att annan enhet väljs för lokal panel
ImageIndexShortCutp�    TActionToolBar2ActionTagCategoryViewCaption   Verktygsfält snabb&tangenterHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för snabbtangenter  TActionCommanderMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHint   Dölj/visa meny  TActionCommanderSessionBandActionTagCategoryViewCaptionSessio&nsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sessioner  TActionCommanderPreferencesBandActionTagCategoryViewCaption   InställningsknapparHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för inställningar  TActionCommanderSortBandActionTagCategoryViewCaptionS&orteringsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sortering  TActionCommanderUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfält för uppdatering  TActionCommanderTransferBandActionTagCategoryViewCaption   ÖverföringsinställningarHelpKeywordui_toolbarsHint9   Dölj/visa verktygsfält för överföringsinställningar  TActionCommanderCommandsBandActionTagCategoryViewCaption&KommandoknapparHelpKeywordui_toolbarsHint)   Visa/dölj verktygsfältet för kommandon  TAction!CommanderCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionCommanderLocalHistoryBandActionTagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för lokal historik  TAction"CommanderLocalNavigationBandActionTagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint0   Dölj/visa verktygsfältet för lokal navigering  TActionCommanderLocalFileBandActionTagCategoryViewCaption&FilknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfältet för lokala filer  TAction!CommanderLocalSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint6   Dölj/visa verktygsfält för lokala markeringsknappar  TAction CommanderRemoteHistoryBandActionTagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet fjärrhistorik  TAction#CommanderRemoteNavigationBandActionTagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint0   Dölj/visa verktygsfältet för fjärrnavigering  TActionCommanderRemoteFileBandActionTagCategoryViewCaption&FilknapparHelpKeywordui_toolbarsHint+   Dölj/visa verktygsfältet för fjärrfiler  TAction"CommanderRemoteSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint7   Visa/dölj verktygsfältet för fjärrmarkeringsknappar  TActionLocalStatusBarActionTagCategoryViewCaption   Statusf&ältHint*   Dölj/visa den lokala panelens statusfält  TActionRemoteStatusBarActionTagCategoryViewCaption   Statusf&ältHint%   Dölj/visa fjärrpanelens statusfält  TActionLocalSortByNameActionTag	CategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint8Sortera efter namn|Sortera den lokala panelen efter namn
ImageIndexShortCutr@  TActionLocalSortByExtActionTag	CategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintF   Sortera efter filändelse|Sortera den lokala panelen efter filändelse
ImageIndex ShortCuts@  TActionLocalSortBySizeActionTag	CategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHintASortera efter storlek|Sortera den lokala panelen efter filstorlek
ImageIndex#ShortCutu@  TActionLocalSortByAttrActionTag	CategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHint@Sortera efter attribut|Sortera den lokala panelen efter attribut
ImageIndex$ShortCutv@  TActionLocalSortByTypeActionTag	CategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint<Sortera efter filtyp|Sortera den lokala panelen efter filtyp
ImageIndex"  TActionLocalSortByChangedActionTag	CategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintM   Sortera efter senast &ändrad|Sortera den lokala panelen efter senast ändrad
ImageIndex!ShortCutt@  TActionRemoteSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintW   Stigande/fallande|Växla sortering mellan stigande och fallande ordning i fjärrpanelen
ImageIndex%  TActionRemoteSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint3   Sortera efter namn|Sortera fjärrpanelen efter namn
ImageIndexShortCutr@  TActionRemoteSortByExtActionTagCategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintA   Sortera efter filändelse|Sortera fjärrpanelen efter filändelse
ImageIndex ShortCuts@  TActionRemoteSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint<   Sortera efter storlek|Sortera fjärrpanelen efter filstorlek
ImageIndex#ShortCutu@  TActionRemoteSortByRightsActionTagCategorySortCaption   Efter &filrättigheterHelpKeywordui_file_panel#sorting_filesHintI   Sortera efter filrättigheter|Sortera fjärrpanelen efter filrättigheter
ImageIndex$ShortCutv@  TActionRemoteSortByChangedActionTagCategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintH   Sortera efter senast &ändrad|Sortera fjärrpanelen efter senast ändrad
ImageIndex!ShortCutt@  TActionRemoteSortByOwnerActionTagCategorySortCaption   Efter ä&gareHelpKeywordui_file_panel#sorting_filesHint:   Sortera efter ägare|Sortera fjärrpanelen efter filägare
ImageIndex&ShortCutw@  TActionRemoteSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHint8   Sortera efter grupp|Sortera fjärrpanelen efter filgrupp
ImageIndex'ShortCutx@  TActionRemoteSortByTypeActionTagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint7   Sortera efter filtyp|Sortera fjärrkatalog efter filtyp
ImageIndex"  TActionCurrentSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintW   Stigande/fallande|Växla sortering mellan stigande och fallande ordning i aktuell panel
ImageIndex%  TActionCurrentSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint3Sortera efter namn|Sortera aktuell panel efter namn
ImageIndexShortCutr@  TActionCurrentSortByExtActionTagCategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintA   Sortera efter filändelse|Sortera aktuell panel efter filändelse
ImageIndex ShortCuts@  TActionCurrentSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint<Sortera efter storlek|Sortera aktuell panel efter filstorlek
ImageIndex#ShortCutu@  TActionCurrentSortByTypeActionTagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHintLSortera efter filtyp|Sortera aktuell panel efter filtyp (endast lokal panel)
ImageIndex"  TActionCurrentSortByRightsActionTagCategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHintK   Sortera efter attribut|Sortera aktuell panel efter attribut/filrättigheter
ImageIndex$ShortCutv@  TActionCurrentSortByChangedActionTagCategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintH   Sortera efter senast &ändrad|Sortera aktuell panel efter senast ändrad
ImageIndex!ShortCutt@  TActionCurrentSortByOwnerActionTagCategorySortCaption   Efter ä&gareHelpKeywordui_file_panel#sorting_filesHintO   Sortera efter ägare|Sortera aktuell panel efter filägare (endast fjärrpanel)
ImageIndex&ShortCutw@  TActionCurrentSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHintM   Sortera efter grupp|Sortera fjärrpanelen efter filgrupp (endast fjärrpanel)
ImageIndex'ShortCutx@  TActionSortColumnAscendingActionTagCategorySortCaptionSortera stig&andeHelpKeywordui_file_panel#sorting_filesHint(Sortera filer stigande efter vald kolumn
ImageIndex)  TActionSortColumnDescendingActionTagCategorySortCaptionSortera fallan&deHelpKeywordui_file_panel#sorting_filesHint(Sortera filer fallande efter vald kolumn
ImageIndex(  TActionHomepageActionTagCategoryHelpCaptionProdukt&hemsidaHint9   Öppnar webbläsaren och går till applikationens hemsida
ImageIndex*  TActionHistoryPageActionTagCategoryHelpCaption&VersionshistorikHintO   Öppnar webbläsaren och går till webbsida med applikationens versionshistorik  TActionSaveCurrentSessionAction2TagCategorySessionCaption&Spara session som webbplats...HelpKeywordtask_connections#savingHint?Spara session som webbplats|Spara aktuell session som webbplats
ImageIndex+  TActionShowHideRemoteNameColumnActionTagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint5   Visa/dölj namn|Visa/dölj namnkolumn i fjärrpanelen
ImageIndex,  TActionShowHideRemoteExtColumnActionTagCategoryColumnsCaption   &FiländelseHelpKeywordui_file_panel#selecting_columnsHintC   Visa/dölj filändelse|Visa/dölj filändelsekolumn i fjärrpanelen
ImageIndex-  TActionShowHideRemoteSizeColumnActionTagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHint?   Visa/dölj storlek|Visa/dölj filstorlekskolumn i fjärrpanelen
ImageIndex/  TAction!ShowHideRemoteChangedColumnActionTagCategoryColumnsCaption   Se&nast ändradHelpKeywordui_file_panel#selecting_columnsHintJ   Visa/dölj senast ändrad|Visa/dölj senast ändrad-kolumn i fjärrpanelen
ImageIndex0  TAction ShowHideRemoteRightsColumnActionTagCategoryColumnsCaption   Fil&rättigheterHelpKeywordui_file_panel#selecting_columnsHintJ   Visa/dölj filrättigheter|Visa/dölj filrättighetskolumn i fjärrpanelen
ImageIndex1  TActionShowHideRemoteOwnerColumnActionTagCategoryColumnsCaption   &ÄgareHelpKeywordui_file_panel#selecting_columnsHint8   Visa/dölj ägare|Visa/dölj ägarkolumn i fjärrpanelen
ImageIndex2  TActionShowHideRemoteGroupColumnActionTagCategoryColumnsCaption&GruppHelpKeywordui_file_panel#selecting_columnsHint7   Visa/dölj grupp|Visa/dölj gruppkolumn i fjärrpanelen
ImageIndex3  TAction$ShowHideRemoteLinkTargetColumnActionTagCategoryColumnsCaption
   &LänkmålHelpKeywordui_file_panel#selecting_columnsHint@   Visa/dölj länkmål|Visa/dölj länkmålskolumn i fjärrpanelen
ImageIndexR  TActionShowHideRemoteTypeColumnActionTagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint:   Visa/dölj filtyp|Visa/dölj filtypskolumn i fjärrpanelen
ImageIndex.  TActionShowHideLocalNameColumnActionTagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint:   Visa/dölj namn|Visa/dölj namnkolumn i den lokala panelen
ImageIndex,  TActionShowHideLocalExtColumnActionTagCategoryColumnsCaption   &FiländelseHelpKeywordui_file_panel#selecting_columnsHintH   Visa/dölj filändelse|Visa/dölj filändelsekolumn i den lokala panelen
ImageIndex-  TActionShowHideLocalTypeColumnActionTagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint?   Visa/dölj filtyp|Visa/dölj filtypskolumn i den lokala panelen
ImageIndex.  TActionShowHideLocalSizeColumnActionTagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHintD   Visa/dölj storlek|Visa/dölj filstorlekskolumn i den lokala panelen
ImageIndex/  TAction ShowHideLocalChangedColumnActionTagCategoryColumnsCaption   Senast &ändradHelpKeywordui_file_panel#selecting_columnsHintO   Visa/dölj senast ändrad|Visa/dölj senast ändrad-kolumn i den lokala panelen
ImageIndex0  TActionShowHideLocalAttrColumnActionTagCategoryColumnsCaption	&AttributHelpKeywordui_file_panel#selecting_columnsHintB   Visa/dölj attribut|Visa/dölj attributkolumn i den lokala panelen
ImageIndex1  TActionCompareDirectoriesActionTagCategoryCommandCaption   &Jämför katalogerHelpKeywordtask_compare_directoriesHintH   Jämför kataloger|Markerar skillnader mellan lokal- och fjärrkatalogen
ImageIndex4ShortCutq   TActionSynchronizeActionTagCategoryCommandCaption!   &Håll fjärrkatalogen uppdateradHelpKeywordtask_keep_up_to_dateHintA   Håll fjärrkatalogen uppdaterad|Håll fjärrkatalogen uppdaterad
ImageIndex5ShortCutU@  TActionForumPageActionTagCategoryHelpCaption&SupportforumHint=   Öppnar webbläsaren och gå till webbsida med supportforumet  TActionLocalAddBookmarkActionTag	CategoryLocal DirectoryCaption   &Lägg till bokmärkenHelpKeywordtask_navigate#bookmarksHintD   Lägg till bokmärken|Lägg till aktuell lokal katalog som bokmärke
ImageIndex6ShortCutB@  TActionRemoteAddBookmarkActionTagCategoryRemote DirectoryCaption   &Lägg till bokmärkenHelpKeywordtask_navigate#bookmarksHintD   Lägg till bokmärken|Lägg till aktuell fjärrkatalog som bokmärke
ImageIndex6ShortCutB@  TActionConsoleActionTagCategoryCommandCaption   Öppna &terminalfönsterHelpKeyword
ui_consoleHint�   Öppna terminalfönster|Öppnar terminalfönster som tillåter körande av godtyckligt extrakommando (med undantag av de som kräver användarinput)
ImageIndex7ShortCutT`  TActionPuttyActionTagCategoryCommandCaption   Öppna session i &PuTTYHelpKeywordintegration_putty#open_puttyHintZ   Öppna session i PuTTY|Starta PuTTY SSH-terminalprogram och öppna aktuell session med den
ImageIndex@ShortCutP@  TActionLocalExploreDirectoryActionTagCategoryLocal DirectoryCaption&Utforska katalogHint+   Öppnar utforskaren i aktuell lokal katalog
ImageIndex8ShortCutE�    TActionCurrentOpenActionTagCategoryFocused OperationCaption   &ÖppnaHelpKeyword	task_editHintQ   Öppna dokument|Öppnar valt dokument med program som filtypen är associerad med
ImageIndex:  TActionSynchronizeBrowsingActionTagCategoryCommand	AutoCheck	Caption   Synkronisera &bläddringHelpKeyword"task_navigate#synchronize_browsingHintJ   Synkronisera bläddring|Synkronisera lokal och fjärrkatalogens bläddring
ImageIndex;ShortCutB�    TActionCurrentAddEditLinkActionTagCategorySelected OperationCaption   Lägg till/redigera &länk...HelpKeyword	task_linkHintZ   Lägg till/redigera länk|Lägger till ny länk/genväg eller redigerar vald länk/genväg
ImageIndex<  TActionCurrentAddEditLinkContextActionTagCategorySelected OperationCaption   Redigera &länk...HelpKeyword	task_linkHint*   Redigera länk|Redigera vald länk/genväg
ImageIndex<  TActionCloseApplicationActionTagCategoryCommandCaption&AvslutaHintG   Avsluta applikation|Avsluta öppnade sessioner och stäng applikationen  TActionOpenedSessionsActionTagCategorySessionCaption   &Öppna sessionerHelpKeywordtask_connections#switchHint0   Välj session|Välj öppnad session att aktivera
ImageIndex>  TActionDuplicateSessionActionTagCategorySessionCaption&Dubblera sessionHelpKeywordtask_connectionsHintf   Dubblera session|Öppnar samma session igen (håll nere SHIFT för att öppna den i ett nytt fönster)
ImageIndex[  TActionNewLinkActionTagCategoryCommandCaption	   &Länk...HelpKeyword	task_linkHint"   Skapa länk|Skapa ny länk/genväg
ImageIndex<  TActionCustomCommandsFileActionTagCategoryCommandCaptionFiler &anpassade kommandonHelpKeywordcustom_commandHint%   Kör anpassade kommandon på vald fil  TActionCustomCommandsNonFileActionTagCategoryCommandCaptionStatiska &anpassade kommandonHelpKeywordcustom_commandHint4   Kör anpassade kommandon som inte fungerar på filer  TActionCustomCommandsCustomizeActionTagCategoryCommandCaption&Anpassa...HelpKeywordui_pref_commandsHintAnpassa egna kommandon
ImageIndex  TActionCustomCommandsEnterActionTagCategoryCommandCaption   Lä&gg in...HelpKeyword(custom_command#executing_and_configuringHint#   Lägg in egna kommandon för ad hoc
ImageIndexZ  TAction CustomCommandsEnterFocusedActionTagCategoryCommandCaption   Lä&gg in...HelpKeyword(custom_command#executing_and_configuringHint#   Lägg in egna kommandon för ad hoc
ImageIndexZ  TActionCheckForUpdatesActionTagCategoryHelpCaption   Sök efter &uppdateringarHelpKeywordupdatesHint0   Frågar applikationens webbsida om uppdateringar
ImageIndex?  TActionDonatePageActionTagCategoryHelpCaption&DoneraHintG   Öppnar webbläsaren och går till programmets webbsida för donationer  TActionCustomCommandsLastActionTagCategoryCommandCaptionCustomCommandsLastActionHelpKeyword(custom_command#executing_and_configuring  TActionCustomCommandsLastFocusedActionTagCategoryCommandCaptionCustomCommandsLastFocusedActionHelpKeyword(custom_command#executing_and_configuring  TActionFileSystemInfoActionTagCategoryCommandCaption&Server/protokollinformationHelpKeyword	ui_fsinfoHint Visa server/protokollinformation
ImageIndex  TActionClearCachesActionTagCategoryCommandCaption&Rensa cacheHelpKeyworddirectory_cacheHint1   Rensa cache för kataloglistning och katalogbyten  TActionFullSynchronizeActionTagCategoryCommandCaption&Synkronisera...HelpKeywordtask_synchronize_fullHint,   Synkronisera lokal katalog med fjärrkatalog
ImageIndexBShortCutS@  TActionRemoteMoveToFocusedActionTagCategoryRemote Focused OperationCaption&Flytta till...HelpKeywordtask_move_duplicate#moveHint0   Flytta|Flytta markerade filer till fjärrkatalog
ImageIndexd  TActionShowHiddenFilesActionTagCategoryViewCaption   Visa/dölj &dolda filerHelpKeywordui_file_panel#hidden_filesHint)   Växla visning av dolda filer i panel(er)ShortCutH�    TActionFormatSizeBytesNoneActionTagCategoryViewCaption&ByteHelpKeywordui_pref_panels#commonHintVisa filstorlekar i byte  TActionLocalPathToClipboardActionTagCategoryLocal DirectoryCaption   Kopiera s&ökväg till urklippHelpKeywordfilenames#cwdHint+   Kopiera aktuell lokal sökväg till urklipp  TActionRemotePathToClipboardActionTagCategoryRemote DirectoryCaption   Kopiera s&ökväg till urklippHelpKeywordfilenames#cwdHint+   Kopiera aktuell fjärrsökväg till urklipp  TActionFileListToCommandLineActionTagCategorySelected OperationCaptionIn&foga till kommandoradHelpKeywordfilenames#command_lineHint/Infoga markerade filers namn till kommandoradenShortCut@  TActionFileListToClipboardActionTagCategorySelected OperationCaption&Kopiera till urklippHelpKeywordfilenames#file_nameHint*Kopiera markerade filers namn till urklippShortCutC`  TActionFullFileListToClipboardActionTagCategorySelected OperationCaption,   Kopiera till urklipp (inklusive s&ökvägar)HelpKeywordfilenames#file_nameHint=   Kopiera markerade filers namn inklusive sökväg till urklippShortCutC�    TActionQueueGoToActionTagCategoryQueueCaption	   &Gå tillHelpKeywordui_queue#manageHint   Gå till överföringskölistan
ImageIndexJShortCutQ@  TActionQueueItemUpActionTagCategoryQueueCaptionFlytta &uppHelpKeywordui_queue#manageHint2   Flytta upp vald köpost för att utföras tidigare
ImageIndexH  TActionQueueItemDownActionTagCategoryQueueCaptionFlytta &nerHelpKeywordui_queue#manageHint0   Flytta ner vald köpost för att utföras senare
ImageIndexI  TActionQueueToggleShowActionTagCategoryQueueCaption   &KöHint   Visa/dölj kölista
ImageIndexJ  TActionQueueShowActionTagCategoryQueueCaptionVi&saHelpKeywordui_queueHint   Visa kölista  TActionQueueHideWhenEmptyActionTagCategoryQueueCaption   Dölj ifall &tomHelpKeywordui_queueHint    Dölj kölistan när den är tom  TActionQueueHideActionTagCategoryQueueCaption   &DöljHelpKeywordui_queueHint   Dölj kölista  TActionQueueToolbarActionTagCategoryQueueCaption   &VerktygsfältHint@   Dölj/visa verktygsfältet för kölistan (på kölistans panel)  TActionQueueFileListActionTagCategoryQueueCaption	&FillistaHint#   Dölj/visa fullständig köfillista  TActionQueuePreferencesActionTagCategoryQueueCaptionA&npassa...HelpKeywordui_pref_backgroundHint   Anpassa kölista
ImageIndex  TActionPasteAction2TagCategoryCommandCaptionK&listra inHelpKeyword	clipboardHint�   Klistra in filer från urklipp till aktuell katalog i aktiv panel; eller öppnar sökväg från urklipp i aktiv panel; eller öppnar sessions-URL från urklipp
ImageIndexKShortCutV@  TActionNewFileActionTagCategoryCommandCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TActionEditorListCustomizeActionTagCategoryCommandCaption&Konfigurera...HelpKeywordui_pref_editorHint   Skräddarsy editorer
ImageIndex  TActionRemoteCopyToFocusedActionTagCategoryRemote Focused OperationCaption&Dubblera...HelpKeywordtask_move_duplicate#duplicateHint3   Dubblera|Dubbleras valda filer till fjärrkatalogen
ImageIndexN  TActionRemoteCopyToActionTagCategoryRemote Selected OperationCaption&Dubblera...HelpKeywordtask_move_duplicate#duplicateHint2   Dubblera|Dubblera valda filer till fjärrkatalogen
ImageIndexN  TActionFileGenerateUrlAction2TagCategorySelected OperationCaptionSkapa fil-&URL...HelpKeywordui_generateurlHint   Skapa URL:er för valda filer  TActionTableOfContentsActionTagCategoryHelpCaption
   I&nnehållHintI   Öppnar webbläsare och går till dokumentationens innehållsförteckning
ImageIndexOShortCutp  TActionFileListFromClipboardActionTagCategorySelected OperationCaption&Transfer Files in ClipboardHelpKeyword	clipboardHint+Transfer files whose names are in clipboard  TActionLocalCopyActionTag	CategoryLocal Selected OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionCurrentDeleteAlternativeActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort valda filer
ImageIndex  TActionCurrentEditWithActionTagCategorySelected OperationCaptionRedigera &med...HelpKeyword	task_editHint9Redigera med|Redigera valda filer med editorn som ni valt  TActionDownloadPageActionTagCategoryHelpCaption
Ladda &nerHintA   Öppnar webbläsare och går till applikationens nerladdningssida  TActionUpdatesPreferencesActionTagCategoryHelpCaptionKonfi&gurera...HelpKeywordui_pref_updatesHintC   Konfigurera automatisk kontroll av uppdateringar för applikationen
ImageIndex  TActionFormatSizeBytesKilobytesActionTagCategoryViewCaption	&KilobyteHelpKeywordui_pref_panels#commonHintVisa filstorlekar i kilobyte  TActionFormatSizeBytesShortActionTagCategoryViewCaption&Kort formatHelpKeywordui_pref_panels#commonHintVisa filstorlekar i kort format  TActionPresetsPreferencesActionTagCategoryViewCaption&Konfigurera...HelpKeywordui_pref_transferHint2   Konfigurera förinställningar för överföringar
ImageIndex  TActionLockToolbarsActionTagCategoryViewCaption   &Lås verktygsfältHelpKeywordui_toolbarsHint3   Hindra flyttning och dockning av alla verktygsfält  TActionSelectiveToolbarTextActionTagCategoryViewCaption&Visa valbara textetiketterHelpKeywordui_toolbarsHintD   Visa textetiketter på utvalda viktiga kommandon på verktygsfältet  TActionCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionColorMenuActionTagCategoryViewCaption   F&ärgHelpKeywordtask_connections#session_colorHint    Ändra färg på aktuell session  TActionAutoReadDirectoryAfterOpActionTagCategoryViewCaptionLadda auto&matisk om katalogHint=   Ändra automatisk omladdning av fjärrkatalog efter operationShortCutR�    TActionQueueItemPauseActionTagCategoryQueueCaption&PausaHelpKeywordui_queue#manageHint   Pausa vald köpost
ImageIndexS  TActionQueueItemResumeActionTagCategoryQueueCaption   &ÅterupptaHelpKeywordui_queue#manageHint   Återuppta vald pausad köpost
ImageIndexF  TActionQueuePauseAllActionTagCategoryQueueCaption&Pausa allaHelpKeywordui_queue#manageHint   Pausa alla köposter som körs
ImageIndexT  TActionQueueResumeAllActionTagCategoryQueueCaption   &Återuppta allaHelpKeywordui_queue#manageHint!   Återuppta alla pausade köposter
ImageIndexU  TActionQueueDeleteAllDoneActionTagCategoryQueueCaption   Ta bort alla &slutfördaHelpKeywordui_queue#manageHint!   Ta bort alla slutförda köposter
ImageIndexc  TActionQueueEnableActionTagCategoryQueueCaption   &ProcessköHelpKeywordui_queue#manageHints   Aktivera köbehandling|Aktivera köbehandling (väntande köposter startar inte, när köbehandling är inaktiverad
ImageIndex`ShortCutQ`  TActionQueueDisconnectOnceEmptyAction2TagCategoryQueueCaption   &Koppla ifrån sessionHelpKeywordui_queueHint'   Koppla ifrån session när kön är tom
ImageIndexW  TActionRestoreSelectionActionTagCategory	SelectionCaption   &Återställ markeringHelpKeywordui_file_panel#selecting_filesHint"   Återställ föregående markering
ImageIndexV  TActionLocalSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint'Markera|Markera lokala filer efter mask
ImageIndex  TActionLocalUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint+Avmarkera|Avmarkera lokala filer efter mask
ImageIndex  TActionLocalSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla lokala filer
ImageIndex  TActionCurrentEditFocusedActionTagCategoryFocused OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera valda filer
ImageIndex9  TActionCurrentEditWithFocusedActionTagCategoryFocused OperationCaptionRedigera &med...HelpKeyword	task_editHint9Redigera med|Redigera valda filer med editorn som ni valt  TActionNewDirActionTagCategoryCommandCaptionKatalo&g...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionQueueShutDownOnceEmptyAction2TagCategoryQueueCaption   Stäng av datornHelpKeywordui_queueHint"   Stäng av datorn när kön är tom
ImageIndex]  TActionQueueSuspendOnceEmptyAction2TagCategoryQueueCaption   Försätt datorn i vilolägeHelpKeywordui_queueHint.   Försätt datorn i viloläge när kön är tom
ImageIndexi  TActionQueueIdleOnceEmptyActionTagCategoryQueueCaption   &Förbli inaktivChecked	HelpKeywordui_queueHint!   Förbli inaktiv när kön är tom
ImageIndex^  TActionQueueCycleOnceEmptyActionTagCategoryQueueCaption   &Tom köHelpKeywordui_queueHint1   Ändra åtgärd som ska utföras då kön är tom
ImageIndex^  TTBEditActionQueueItemSpeedActionTagCategoryQueueHelpKeywordui_queue#manageHint)   Ändra hastighetsgräns för vald köpost
ImageIndexmEditCaption
&Hastighet  TActionQueueDeleteAllActionTagCategoryQueueCaption&Avbryt allaHelpKeywordui_queue#manageHint   Ta bort alla köposter
ImageIndexj  TActionLocalFilterActionTag	CategoryLocal DirectoryCaption&Filtrera...HelpKeywordui_file_panel#filteringHintFiltrera|Filtrera visade filer
ImageIndex\ShortCutF�    TActionRemoteFilterActionTagCategoryRemote DirectoryCaption
&Filter...HelpKeywordui_file_panel#filteringHintFilter|Filtrera visade filer
ImageIndex\ShortCutF�    TActionRemoteFindFilesActionTagCategoryRemote DirectoryCaption   Sö&k filer..HelpKeyword	task_findHint#   Sök filer|Sök filer och kataloger
ImageIndex_  TActionCurrentEditInternalActionTagCategorySelected OperationCaption&Intern editorHelpKeyword	task_editHint8Redigera (intern)|Redigera valda filer med intern editor  TActionSaveWorkspaceActionTagCategorySessionCaptionSpara arbets&yta...HelpKeyword	workspaceHintSpara arbetsyta|Spara arbetsyta
ImageIndexf  TActionLocalRenameActionTagCategoryLocal Selected OperationCaption	&Byt namnHelpKeywordtask_renameHint$   Byt namn|Byt namn på vald lokal fil
ImageIndex  TActionLocalEditActionTagCategoryLocal Selected OperationCaption	&RedigeraHelpKeyword	task_editHint$Redigera|Redigera valda lokala filer
ImageIndex9  TActionLocalMoveActionTag	CategoryLocal Selected OperationCaption   Överför och ta &bort...HelpKeywordtask_uploadHint]   Överför och ta bort|Överför valda lokala filer till fjärrkatalogen och tar bort original
ImageIndexb  TActionLocalCreateDirAction2TagCategoryLocal Selected OperationCaptionKatalo&g...HelpKeywordtask_create_directoryHint$Skapa katalog|Skapa ny lokal katalog
ImageIndex  TActionLocalDeleteActionTagCategoryLocal Selected OperationCaption&Ta bortHelpKeywordtask_deleteHint"Ta bort|Ta bort valda lokala filer
ImageIndex  TActionLocalPropertiesActionTagCategoryLocal Selected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint9   Egenskaper|Visa/ändra egenskaper för valda lokala filer
ImageIndex  TActionLocalAddEditLinkAction2TagCategoryLocal Selected OperationCaption   &Genväg...HelpKeyword	task_linkHint\   Lägg till/redigera genväg|Lägg till en ny lokal genväg eller redigera vald lokal genväg
ImageIndex<  TActionRemoteRenameActionTagCategoryRemote Selected OperationCaption	&Byt namnHelpKeywordtask_renameHint$   Byt namn|Byt namn på vald fjärrfil
ImageIndex  TActionRemoteEditActionTagCategoryRemote Selected OperationCaption	&RedigeraHelpKeyword	task_editHint#   Redigera|Redigera valda fjärrfiler
ImageIndex9  TActionRemoteMoveActionTagCategoryRemote Selected OperationCaptionLadda ner och &ta bortHelpKeywordtask_downloadHintY   Ladda ner och ta bort|Ladda ner valda fjärrfiler till lokal katalog och ta bort original
ImageIndexa  TActionRemoteCreateDirAction2TagCategoryRemote Selected OperationCaptionKatalo&g...HelpKeywordtask_create_directoryHint$   Skapa katalog|Skapa ny fjärrkatalog
ImageIndex  TActionRemoteDeleteActionTagCategoryRemote Selected OperationCaption&Ta bortHelpKeywordtask_deleteHint!   Ta bort|Ta bort valda fjärrfiler
ImageIndex  TActionRemotePropertiesActionTagCategoryRemote Selected OperationCaption&EgenskaperHelpKeywordtask_propertiesHintZ   Egenskaper|Visa/ändra rättigheter, ägarskap och andra egenskaper för valda fjärrfiler
ImageIndex  TActionRemoteAddEditLinkAction2TagCategoryRemote Selected OperationCaption	   &Länk...HelpKeyword	task_linkHintQ   Lägg till/ändra länk|Lägg till ny fjärrlänk eller redigera vald fjärrlänk
ImageIndex<  TActionRemoteSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint&   Markera|Markera fjärrfiler efter mask
ImageIndex  TActionRemoteUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint*   Avmarkera|Avmarkera fjärrfiler efter mask
ImageIndex  TActionRemoteSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHint   Markera alla fjärrfiler
ImageIndex  TActionLocalMoveFocusedActionTagCategoryLocal Focused OperationCaption   Överför och &ta bort...HelpKeywordtask_uploadHintZ   Överför och ta bort|Överför valda lokala filer till fjärrkatalog och ta bort original
ImageIndexb  TAction CurrentEditInternalFocusedActionTagCategoryFocused OperationCaption&Intern editorHelpKeyword	task_editHint8Redigera (intern)|Redigera valda filer med intern editor  TActionCurrentSystemMenuFocusedActionTagCategoryFocused OperationCaption&SystemmenyHintn   Visa filsystemets snabbmeny (i egenskaper kan du välja att visa den som standard istället för inbyggd meny)  TActionSessionGenerateUrlAction2TagCategorySessionCaptionSkapa sessions-&URL/kod...HelpKeywordui_generateurlHint/   Skapa URL eller kod för den aktuella sessionen  TActionSelectSameExtActionTagCategory	SelectionCaption$   &Markera filer med samma filtilläggHint:   Markera alla filer med samma filtillägg som fokuserad filShortCutk�    TActionUnselectSameExtActionTagCategory	SelectionCaption&   &Avmarkera filer med samma filtilläggHint<   Avmarkera alla filer med samma filtillägg som fokuserad filShortCutm�    TActionGoToAddressActionTagCategoryCommandCaptionGoToAddressActionSecondaryShortCuts.StringsAlt+D ShortCutL@  TAction
LockActionTagCategorySelected OperationCaption   &LåsHint   Lås markerade filer  TActionUnlockActionTagCategorySelected OperationCaption	   Lås &uppHint   Lås upp markerade filer  TAction
TipsActionTagCategoryHelpCaption
Visa &tipsHelpKeywordui_tipsHint%   Visar tips om hur du använder WinSCP
ImageIndexn  TActionChangePasswordActionTagCategorySessionCaption   Ä&ndra lösenord...HelpKeywordtask_change_passwordHint   Ändra kontolösenord  TActionPrivateKeyUploadActionTagCategorySessionCaption,&Installera den publika nyckeln i servern...HelpKeywordguide_public_keyHint;   Installera den publika nyckeln för autentisering i servern  TActionRemoteNewFileActionTagCategoryRemote Selected OperationCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TActionLocalNewFileActionTagCategoryLocal Selected OperationCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TActionCustomizeToolbarActionTagCategoryViewCaption   &Anpassa verktygsfältetHelpKeywordui_toolbarsHint    Visa/dölj verktygsfältsknappar  TActionRenameSessionActionTagCategorySessionCaption   &Byt namn på sessionHelpKeywordtask_connections#renamingHint<   Byt namn på session|Ändrar namn på den aktuella sessionen  TActionCurrentCopyToClipboardActionTagCategorySelected OperationCaptionK&opieraHelpKeywordclipboard#copyHint-Kopiera|Kopiera de valda filerna till urklipp
ImageIndexoShortCutC@  TActionFileColorsPreferencesActionTagCategoryViewCaption   Fil&färger...HelpKeywordui_pref_file_colorsHint   Konfigurera filfärgsregler  TAction#CurrentCopyToClipboardFocusedActionTagCategoryFocused OperationCaptionK&opieraHelpKeywordclipboard#copyHint-Kopiera|Kopiera de valda filerna till urklipp
ImageIndexoShortCutC@   TTBXPopupMenuExplorerBarPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left� TopP TTBXItemAddress2ActionExplorerAddressBandAction  TTBXItemStandardButtons1ActionExplorerToolbarBandAction  TTBXItemSelectionButtons1ActionExplorerSelectionBandAction  TTBXItemSessionButtons2ActionExplorerSessionBandAction  TTBXItemPreferencesButtons1ActionExplorerPreferencesBandAction  TTBXItemSortButtons3ActionExplorerSortBandAction  TTBXItemTBXItem3ActionExplorerUpdatesBandAction  TTBXItemTBXItem4ActionExplorerTransferBandAction  TTBXItem	TBXItem16Action ExplorerCustomCommandsBandAction  TTBXItemTBXItem7ActionLockToolbarsAction  TTBXItem	TBXItem48ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem4ActionCustomizeToolbarAction  TTBXSeparatorItemN5  TTBXItemSessionsTabsAction2ActionSessionsTabsAction  TTBXItem
StatusBar2ActionStatusBarAction  TTBXSeparatorItemN72  TTBXSubmenuItemQueue7Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow6ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty6ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide5ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN71  TTBXItemToolbar5ActionQueueToolbarAction  TTBXItem	TBXItem85ActionQueueFileListAction  TTBXSeparatorItemN70  TTBXItem
Customize5ActionQueuePreferencesAction   TTBXItemTree4ActionRemoteTreeAction   TTimerSessionIdleTimerEnabledInterval�OnTimerSessionIdleTimerTimerLeft TopP  TTBXPopupMenuCommanderBarPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�Top TTBXItemCommandsButtons2ActionCommanderCommandsBandAction  TTBXItemSessionButtons5ActionCommanderSessionBandAction  TTBXItemPreferencesButtons4ActionCommanderPreferencesBandAction  TTBXItemSortButtons2ActionCommanderSortBandAction  TTBXItemTBXItem2ActionCommanderUpdatesBandAction  TTBXItemTBXItem5ActionCommanderTransferBandAction  TTBXItem	TBXItem15Action!CommanderCustomCommandsBandAction  TTBXItemTBXItem6ActionLockToolbarsAction  TTBXItem	TBXItem46ActionSelectiveToolbarTextAction  TTBXSubmenuItem	TBXItem77ActionCustomizeToolbarAction  TTBXSeparatorItemN26  TTBXItemSessionsTabsAction1ActionSessionsTabsAction  TTBXItemCommandLine2ActionCommandLinePanelAction  TTBXItemCommandsToolbar1ActionToolBar2Action  TTBXItem
StatusBar8ActionStatusBarAction  TTBXSeparatorItemN27  TTBXSubmenuItemLocalPanel1Caption&Lokal panelHelpKeywordui_file_panelHint#   Ändra den lokala panelens utseende TTBXItemHistoryButtons3ActionCommanderLocalHistoryBandAction  TTBXItemNavigationButtons3Action"CommanderLocalNavigationBandAction  TTBXItem	TBXItem40ActionCommanderLocalFileBandAction  TTBXItem	TBXItem43Action!CommanderLocalSelectionBandAction  TTBXSeparatorItemN23  TTBXItemTree7ActionLocalTreeAction  TTBXSeparatorItemN77  TTBXItem
StatusBar6ActionLocalStatusBarAction   TTBXSubmenuItemRemotePanel2Caption   &FjärrpanelHelpKeywordui_file_panelHint   Ändra fjärrpanelens utseende TTBXItemHistoryButtons4Action CommanderRemoteHistoryBandAction  TTBXItemNavigationButtons4Action#CommanderRemoteNavigationBandAction  TTBXItem	TBXItem41ActionCommanderRemoteFileBandAction  TTBXItem	TBXItem42Action"CommanderRemoteSelectionBandAction  TTBXSeparatorItemN25  TTBXItemTree8ActionRemoteTreeAction  TTBXSeparatorItemN78  TTBXItem
StatusBar7ActionRemoteStatusBarAction   TTBXSubmenuItemOptions1Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow5ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty5ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide4ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN69  TTBXItemToolbar4ActionQueueToolbarAction  TTBXItem	TBXItem84ActionQueueFileListAction  TTBXSeparatorItemN68  TTBXItem
Customize4ActionQueuePreferencesAction    TTBXPopupMenuRemotePanelPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left8Top TTBXSubmenuItemTBXSubmenuItem8Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem86ActionRemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem13  TTBXItem	TBXItem87ActionRemoteParentDirAction  TTBXItem	TBXItem88ActionRemoteRootDirAction  TTBXItem	TBXItem89ActionRemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem90ActionRemoteBackAction  TTBXItem	TBXItem91ActionRemoteForwardAction   TTBXItem	TBXItem32ActionRemoteRefreshAction  TTBXItem	TBXItem30ActionRemoteAddBookmarkAction  TTBXItem	TBXItem26ActionRemoteFilterAction  TTBXItemCopyPathtoClipboard1ActionRemotePathToClipboardAction  TTBXSeparatorItemN51  TTBXItemHistoryButtons5Action CommanderRemoteHistoryBandAction  TTBXItemNavigationButtons5Action#CommanderRemoteNavigationBandAction  TTBXItem	TBXItem14ActionCommanderRemoteFileBandAction  TTBXItem	TBXItem45Action"CommanderRemoteSelectionBandAction  TTBXItem	TBXItem37ActionLockToolbarsAction  TTBXItem	TBXItem49ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem9ActionCustomizeToolbarAction  TTBXSeparatorItemN28  TTBXItemTree5ActionRemoteTreeAction  TTBXSeparatorItemN75  TTBXItem
StatusBar9ActionRemoteStatusBarAction   TTBXPopupMenuLocalPanelPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left8TopP TTBXSubmenuItemTBXSubmenuItem10Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem92ActionLocalOpenDirAction  TTBXItem	TBXItem93ActionLocalExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem	TBXItem94ActionLocalParentDirAction  TTBXItem	TBXItem95ActionLocalRootDirAction  TTBXItem	TBXItem96ActionLocalHomeDirAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem97ActionLocalBackAction  TTBXItem	TBXItem98ActionLocalForwardAction   TTBXItem	TBXItem34ActionLocalRefreshAction  TTBXItem	TBXItem27ActionLocalFilterAction  TTBXItem	TBXItem31ActionLocalAddBookmarkAction  TTBXItemCopyPathtoClipboard2ActionLocalPathToClipboardAction  TTBXSeparatorItemN52  TTBXItemHistoryButtons6ActionCommanderLocalHistoryBandAction  TTBXItemNavigationButtons6Action"CommanderLocalNavigationBandAction  TTBXItem	TBXItem39ActionCommanderLocalFileBandAction  TTBXItem	TBXItem44Action!CommanderLocalSelectionBandAction  TTBXItem	TBXItem38ActionLockToolbarsAction  TTBXItem	TBXItem47ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem6ActionCustomizeToolbarAction  TTBXSeparatorItemN29  TTBXItemTree6ActionLocalTreeAction  TTBXSeparatorItemN76  TTBXItemStatusBar10ActionLocalStatusBarAction   TTBXPopupMenuLocalDirViewColumnPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left� TopX TTBXItemSortAscending1ActionSortColumnAscendingAction  TTBXItemSortDescending1ActionSortColumnDescendingAction  TTBXItemLocalSortByExtColumnPopupItemActionLocalSortByExtAction  TTBXItemHidecolumn1ActionHideColumnAction  TTBXSeparatorItemN37  TTBXSubmenuItemLocalFormatSizeBytesPopupItemCaptionVisa &filstorlekar iHelpKeywordui_pref_panels#commonHint$   Välj visningsformat för filstorlek TTBXItem	TBXItem64ActionFormatSizeBytesNoneAction  TTBXItem	TBXItem65ActionFormatSizeBytesKilobytesAction  TTBXItem	TBXItem66ActionFormatSizeBytesShortAction   TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItemShowcolumns3CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint&   Välj kolumner som ska visas i panelen TTBXItemName3ActionShowHideLocalNameColumnAction  TTBXItemSize3ActionShowHideLocalSizeColumnAction  TTBXItemType2ActionShowHideLocalTypeColumnAction  TTBXItemModification3Action ShowHideLocalChangedColumnAction  TTBXItemAttributes3ActionShowHideLocalAttrColumnAction    TTBXPopupMenuRemoteDirViewColumnPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�TopX TTBXItem	MenuItem1ActionSortColumnAscendingAction	RadioItem	  TTBXItem	MenuItem2ActionSortColumnDescendingAction	RadioItem	  TTBXItemRemoteSortByExtColumnPopupItemActionRemoteSortByExtAction  TTBXItemHidecolumn2ActionHideColumnAction  TTBXSeparatorItemN38  TTBXSubmenuItemRemoteFormatSizeBytesPopupItemCaptionVisa &filstorlekar iHelpKeywordui_pref_panels#commonHint$   Välj visningsformat för filstorlek TTBXItem	TBXItem67ActionFormatSizeBytesNoneAction  TTBXItem	TBXItem53ActionFormatSizeBytesKilobytesAction  TTBXItem	TBXItem55ActionFormatSizeBytesShortAction   TTBXSeparatorItemTBXSeparatorItem7  TTBXSubmenuItemShowcolumns4CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint&   Välj kolumner som ska visas i panelen TTBXItemName4ActionShowHideRemoteNameColumnAction  TTBXItemSize4ActionShowHideRemoteSizeColumnAction  TTBXItemTBXItem8ActionShowHideRemoteTypeColumnAction  TTBXItemModification4Action!ShowHideRemoteChangedColumnAction  TTBXItemPermissions1Action ShowHideRemoteRightsColumnAction  TTBXItemOwner2ActionShowHideRemoteOwnerColumnAction  TTBXItemGroup2ActionShowHideRemoteGroupColumnAction  TTBXItemTBXItem1Action$ShowHideRemoteLinkTargetColumnAction    TTBXPopupMenu
QueuePopupImagesGlyphsModule.ExplorerImagesOnPopupQueuePopupPopupOptionstboShowHint Left�Top�  TTBXItem
ShowQuery1ActionQueueItemQueryAction  TTBXItem
ShowError1ActionQueueItemErrorAction  TTBXItemShowPrompt1ActionQueueItemPromptAction  TTBXSeparatorItemN53  TTBXItemExecuteNow1ActionQueueItemExecuteAction  TTBXItemTBXItem9ActionQueueItemPauseAction  TTBXItem	TBXItem10ActionQueueItemResumeAction  TTBXItemDelete4ActionQueueItemDeleteAction  TTBXComboBoxItemQueuePopupSpeedComboBoxItemActionQueueItemSpeedAction	ShowImage	OnAdjustImageIndex+QueuePopupSpeedComboBoxItemAdjustImageIndex  TTBXSeparatorItemN54  TTBXItemMoveUp1ActionQueueItemUpAction  TTBXItem	MoveDown1ActionQueueItemDownAction  TTBXSeparatorItemN67  TTBXItemQueueEnableItemActionQueueEnableAction  TTBXSubmenuItemTBXSubmenuItem1Caption&AllaHelpKeywordui_queue#manageHint&   Administrationskommandon för kömassa TTBXItem	TBXItem11ActionQueuePauseAllAction  TTBXItem	TBXItem12ActionQueueResumeAllAction  TTBXItem
TBXItem142ActionQueueDeleteAllAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem51ActionQueueDeleteAllDoneAction   TTBXSubmenuItemTBXSubmenuItem3ActionQueueCycleOnceEmptyActionDropdownCombo	 TTBXItem	TBXItem28ActionQueueIdleOnceEmptyAction	RadioItem	  TTBXItem	TBXItem13ActionQueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem	TBXItem68ActionQueueSuspendOnceEmptyAction2	RadioItem	  TTBXItem	TBXItem29ActionQueueShutDownOnceEmptyAction2	RadioItem	   TTBXSubmenuItemQueue2Caption&AlternativHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow4ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty4ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide3ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN66  TTBXItemToolbar3ActionQueueToolbarAction  TTBXItem	TBXItem83ActionQueueFileListAction  TTBXSeparatorItemN65  TTBXItem
Customize3ActionQueuePreferencesAction    TTBXPopupMenuRemoteDirViewPopup	AutoPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint LefthTop� TTBXSubmenuItemGoTo4Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemOpenDirectoryBookmark3ActionRemoteOpenDirAction  TTBXSeparatorItemN81  TTBXItemParentDirectory4ActionRemoteParentDirAction  TTBXItemRootDirectory4ActionRemoteRootDirAction  TTBXItemHomeDirectory4ActionRemoteHomeDirAction  TTBXSeparatorItemN80  TTBXItemBack4ActionRemoteBackAction  TTBXItemForward4ActionRemoteForwardAction   TTBXItemRefresh4ActionRemoteRefreshAction  TTBXItemAddToBookmarks4ActionRemoteAddBookmarkAction  TTBXItem	TBXItem35ActionRemoteFilterAction  TTBXItemCopyPathtoClipboard6ActionRemotePathToClipboardAction  TTBXSeparatorItemN79  TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135ActionNewFileAction  TTBXItem
TBXItem136ActionNewDirAction  TTBXItem
TBXItem209ActionNewLinkAction   TTBXItem	TBXItem75ActionPasteAction2  TTBXSubmenuItem$RemoteDirViewPopupCustomCommandsMenuActionCustomCommandsNonFileAction   TTBXPopupMenuLocalDirViewPopup	AutoPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�Top� TTBXSubmenuItemGoTo5Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemOpenDirectoryBookmark4ActionLocalOpenDirAction  TTBXItemExploreDirectory2ActionLocalExploreDirectoryAction  TTBXSeparatorItemN84  TTBXItemParentDirectory5ActionLocalParentDirAction  TTBXItemRootDirectory5ActionLocalRootDirAction  TTBXItemHomeDirectory5ActionLocalHomeDirAction  TTBXSeparatorItemN83  TTBXItemBack5ActionLocalBackAction  TTBXItemForward5ActionLocalForwardAction   TTBXItemRefresh5ActionLocalRefreshAction  TTBXItem	TBXItem36ActionLocalFilterAction  TTBXItemAddToBookmarks5ActionLocalAddBookmarkAction  TTBXItemCopyPathtoClipboard7ActionLocalPathToClipboardAction  TTBXSeparatorItemN82  TTBXSubmenuItemTBXSubmenuItem7Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem	TBXItem70ActionNewFileAction  TTBXItem	TBXItem71ActionNewDirAction   TTBXItem	TBXItem76ActionPasteAction2   TTBXPopupMenuRemoteAddressPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left� Top� TTBXItem	TBXItem33ActionRemoteRefreshAction  TTBXItem	TBXItem24ActionRemoteAddBookmarkAction  TTBXItem	TBXItem25ActionRemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItem	TBXItem17ActionRemoteOpenDirAction  TTBXSubmenuItemTBXSubmenuItem2Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem18ActionRemoteParentDirAction  TTBXItem	TBXItem19ActionRemoteRootDirAction  TTBXItem	TBXItem20ActionRemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem21ActionRemoteBackAction  TTBXItem	TBXItem22ActionRemoteForwardAction    TTBXPopupMenuSessionsPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�Top�  TTBXItem
TBXItem124ActionCloseSessionAction2  TTBXItem	TBXItem79ActionDisconnectSessionAction  TTBXItem	TBXItem80ActionReconnectSessionAction  TTBXItem
TBXItem219ActionDuplicateSessionAction  TTBXItem	TBXItem78ActionRenameSessionAction  TTBXItem
TBXItem125ActionSaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem56ActionFileSystemInfoAction  TTBXItem	TBXItem52ActionSessionGenerateUrlAction2  TTBXSeparatorItemTBXSeparatorItem52  TTBXColorItemColorMenuItemActionColorMenuActionColorclNone  TTBXSeparatorItemTBXSeparatorItem34  TTBXItem
TBXItem123ActionNewSessionAction  TTBXSubmenuItemTBXSubmenuItem23ActionSavedSessionsAction2OptionstboDropdownArrow   TTBXSeparatorItemTBXSeparatorItem35  TTBXItemSessionsTabsAction4ActionSessionsTabsAction   TTBXPopupMenuLocalFilePopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint LeftTopP TTBXItemLocalOpenMenuItemActionCurrentOpenAction  TTBXSubmenuItemLocalEditMenuItemActionCurrentEditFocusedActionDropdownCombo	OnPopupFocusedEditMenuItemPopup  TTBXSubmenuItemLocalCopyMenuItemActionLocalCopyFocusedActionDropdownCombo	 TTBXItem	TBXItem73ActionLocalCopyFocusedNonQueueAction  TTBXItem	TBXItem74ActionLocalCopyFocusedQueueAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem54ActionLocalMoveFocusedAction   TTBXItem	TBXItem57ActionCurrentDeleteFocusedAction  TTBXItem	TBXItem58ActionCurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem81Action#CurrentCopyToClipboardFocusedAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXSubmenuItem LocalFilePopupCustomCommandsMenuActionCustomCommandsFileAction TTBXItem    TTBXSubmenuItemTBXSubmenuItem5Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem59ActionFileListToCommandLineAction  TTBXItem	TBXItem60ActionFileListToClipboardAction  TTBXItem	TBXItem61ActionFullFileListToClipboardAction   TTBXSeparatorItemTBXSeparatorItem4  TTBXItem	TBXItem63ActionCurrentPropertiesFocusedAction  TTBXItem	TBXItem50ActionCurrentSystemMenuFocusedAction       TPF0TOpenDirectoryDialogOpenDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_opendirBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionOpen directoryClientHeightNClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize�N PixelsPerInch`
TextHeight TLabel	EditLabelLeft.TopWidthLHeightCaption   &Öppna katalog:  TImageImageLeftTopWidth Height AutoSize	  THistoryComboBoxLocalDirectoryEditLeft.TopWidthHeightAnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChangeDirectoryEditChangeSaveOn   THistoryComboBoxRemoteDirectoryEditLeft.TopWidth_HeightAnchorsakLeftakTopakRight DropDownCount	MaxLength�TabOrder TextRemoteDirectoryEditOnChangeDirectoryEditChangeSaveOn   TButtonOKBtnLeft� Top,WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top,WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTop8Width�Height� 
ActivePageSessionBookmarksSheetAnchorsakLeftakTopakRightakBottom TabOrderOnChangePageControlChange 	TTabSheetSessionBookmarksSheetTagCaption   Sessionsbokmärken
DesignSizez�   TListBoxSessionBookmarksListTagLeft
Top	WidthHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSessionBookmarkButtonTagLeftTop	WidthSHeightAnchorsakTopakRight Caption   &Lägg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeftTop)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�LeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick   	TTabSheetSharedBookmarksSheetTagCaption   Delade bokmärken
ImageIndex
DesignSizez�   TListBoxSharedBookmarksListTagLeft
Top	WidthHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSharedBookmarkButtonTagLeftTop	WidthSHeightAnchorsakTopakRight Caption   &Lägg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeftTop)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSharedBookmarkButtonTag�LeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeftTopIWidthSHeightAnchorsakTopakRight Caption   &Genväg...TabOrderOnClickShortCutBookmarkButtonClick    TButtonLocalDirectoryBrowseButtonLeft@TopWidthKHeightAnchorsakTopakRight Caption   Blädd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop,WidthyHeightAnchorsakLeftakBottom CaptionP&latsprofiler...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeft@Top,WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TPreferencesDialogPreferencesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption   InställningarClientHeight�ClientWidth!Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize!� PixelsPerInch`
TextHeight TButtonOKButtonLeftTop�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCloseButtonLeftrTop�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPanel	MainPanelLeft Top Width!Height�AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlLeft� Top Width�Height�
ActivePagePreferencesSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetPreferencesSheetTagHelpType	htKeywordHelpKeywordui_pref_environmentCaption   Miljö
ImageIndex
TabVisible
DesignSize��  	TGroupBoxCommonPreferencesGroupLeftTopWidth�Height'AnchorsakLeftakTopakRight Caption   BekräftelserTabOrder 
DesignSize�'  	TCheckBoxSynchronizeSummaryCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption   &SynkroniseringsöversiktTabOrder
OnClickControlChange  	TCheckBoxConfirmOverwritingCheckLeftTopCWidtheHeightAnchorsakLeftakTopakRight Caption   Ö&verskrivning av filerTabOrderOnClickControlChange  	TCheckBoxConfirmDeletingCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption%&Borttagning av filer (rekommenderad)TabOrderOnClickControlChange  	TCheckBoxConfirmClosingSessionCheck2LeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption*   Stäng sessioner när programmet avs&lutasTabOrderOnClickControlChange  	TCheckBoxDDTransferConfirmationCheck2Left Top,WidthUHeightAnchorsakLeftakTopakRight Caption?   D&ra && släpp operationer och klistra in i andra applikationerTabOrderOnClickControlChange  	TCheckBoxContinueOnErrorCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption*   Fortsätt vid &fel (avancerade användare)TabOrderOnClickControlChange  	TCheckBoxConfirmExitOnCompletionCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption.   Avsluta a&pplikationen vid slutförd operationTabOrderOnClickControlChange  	TCheckBoxConfirmResumeCheckLeftTopZWidtheHeightAnchorsakLeftakTopakRight Caption   &Återuppta överföringTabOrderOnClickControlChange  	TCheckBoxConfirmCommandSessionCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption   Öppna separat &skalsessionTabOrder	OnClickControlChange  	TCheckBoxConfirmRecyclingCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption &Flytta filer till papperskorgenTabOrderOnClickControlChange  	TCheckBoxConfirmTransferringCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   &Överföring av filerTabOrder OnClickControlChange  TStaticTextBackgroundConfirmationsLinkLeft TopoWidthYHeight	AlignmenttaRightJustifyAutoSizeCaption/   Ändra bekräftelser av bakgrundsöverföringarTabOrderTabStop	OnClick BackgroundConfirmationsLinkClick   	TGroupBoxNotificationsGroupLeftTop5Width�HeightIAnchorsakLeftakTopakRight CaptionMeddelandenTabOrder
DesignSize�I  TLabelBeepOnFinishAfterTextLeftxTopWidthHeightAnchorsakTopakRight CaptionsShowAccelChar  	TCheckBoxBeepOnFinishCheckLeftTopWidth$HeightAnchorsakLeftakTopakRight Caption=   S&ystemljud när operationen är klar, om den pågår mer änTabOrder OnClickControlChange  TUpDownEditBeepOnFinishAfterEditLeft:TopWidth9Height	AlignmenttaRightJustify	Increment       �@MaxValue      ��@AnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChange  	TCheckBoxBalloonNotificationsCheckLeftTop.WidthlHeightAnchorsakLeftakTopakRight CaptionK   Visa ballong&meddelanden i aktivitetsfältets statusområde (systemfältet)TabOrderOnClickControlChange    	TTabSheetLogSheetTagHelpType	htKeywordHelpKeywordui_pref_loggingCaptionLoggning
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLoggingGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Alternativ för loggningTabOrder 
DesignSize��   TLabelLogMaxSizeCountFilesLabelLeftGTop� WidthHeightCaptionfilerFocusControlLogMaxSizeCountEditShowAccelChar  TLabelLogFileNameLabelLeft(Top.Width.HeightCaption   &Loggsökväg:FocusControlLogFileNameEdit3OnClickControlChange  TFilenameEditLogFileNameEdit3Left(Top>WidthOHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogKinddkSave
DefaultExtlogFilter4Sessionsloggfilar (*.log)|*.log|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för sessionslogg.ClickKey@AnchorsakLeftakTopakRight TabOrderTextLogFileNameEdit3OnChangeControlChange  TPanelLogFilePanelLeft(TopVWidth	HeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder TRadioButtonLogFileAppendButtonLeft TopWidthjHeightCaption   L&ägg tillTabOrder OnClickControlChange  TRadioButtonLogFileOverwriteButtonLeftpTopWidthjHeightCaption   Sk&riv överTabOrderOnClickControlChange   	TComboBoxLogProtocolCombo2Left TopWidthwHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChangeControlChangeItems.Strings	ReduceradNormalDebug 1Debug 2   TStaticTextLogFileNameHintTextLeftTopTWidthoHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  	TCheckBoxEnableLoggingCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption!   Aktivera &sessionslogg på nivå:TabOrder OnClickControlChange  	TCheckBoxLogSensitiveCheckLeft(Top� WidthOHeightAnchorsakLeftakTopakRight Caption/   Logga &lösenord och annan känslig informationTabOrder	OnClickControlChange  	TCheckBoxLogMaxSizeCheckLeft(TopsWidth� HeightAnchorsakLeftakTopakRight Caption$   &Rotera loggfiler efter de har nåttTabOrderOnClickControlChange  	TComboBoxLogMaxSizeComboLeft TopqWidthwHeightAnchorsakTopakRight TabOrderOnChangeControlChangeOnExitLogMaxSizeComboExitItems.Strings1M10M100M1G   	TCheckBoxLogMaxSizeCountCheckLeft@Top� Width� HeightAnchorsakLeftakTopakRight Caption!   &Ta bort gamla loggfiler, behållTabOrderOnClickControlChange  TUpDownEditLogMaxSizeCountEditLeft Top� WidthAHeightMaxValue      ��@MinValue       ��?TabOrderOnChangeControlChange   	TGroupBoxActionsLoggingGroupLeftTop� Width�HeightVAnchorsakLeftakTopakRight CaptionXML-loggTabOrder
DesignSize�V  TFilenameEditActionsLogFileNameEditLeft(Top+WidthOHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogKinddkSave
DefaultExtxmlFilter0XML-loggfiler (*.xml)|*.xml|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för XML-logg.ClickKey@AnchorsakLeftakTopakRight TabOrderTextActionsLogFileNameEditOnChangeControlChange  TStaticTextActionsLogFileNameHintTextLeftTopAWidthoHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   möns&terTabOrderTabStop	  	TCheckBoxEnableActionsLoggingCheckLeftTopWidthgHeightAnchorsakLeftakTopakRight CaptionAktivera &XML-logg till fil:TabOrder OnClickControlChange    	TTabSheetGeneralSheetTagHelpType	htKeywordHelpKeywordui_pref_interfaceCaption   Gränssnitt
ImageIndex
TabVisible
DesignSize��  TLabelInterfaceChangeLabelLeftTopWidth� HeightCaption.   Ändringar kommer att gälla vid nästa start.ShowAccelChar  	TGroupBoxInterfaceGroupLeftTopBWidth�Height� AnchorsakLeftakTopakRightakBottom Caption   AnvändargränssnittTabOrder
DesignSize��   TLabelCommanderDescriptionLabel2Left� TopWidth� HeightsAnchorsakLeftakTopakRight AutoSizeCaption�   - två paneler (vänster för lokal katalog, höger för fjärrkatalog)
- snabbkommandon som i Norton Commander (och andra liknande program som Total Commander, Midnight Commander...)
- dra && släpp till/från båda panelernaWordWrap	OnClickCommanderClick  TLabelExplorerDescriptionLabelLeft� Top� Width� Height>AnchorsakLeftakTopakRight AutoSizeCaptionK   - endast fjärrkatalog
- snabbkommandon som i Utforskaren
- dra && släppWordWrap	OnClickExplorerClick  TImageCommanderInterfacePictureLeft7Top)Width Height AutoSize	OnClickCommanderClick  TImageExplorerInterfacePictureLeft7Top� Width Height AutoSize	OnClickExplorerClick  TRadioButtonCommanderInterfaceButton2LeftTopWidthtHeightCaption
&CommanderChecked	TabOrder TabStop	OnClickControlChange  TRadioButtonExplorerInterfaceButton2LeftTop� WidthoHeightCaption&UtforskareTabOrderOnClickControlChange   	TGroupBox
ThemeGroupLeftTopWidth�Height4AnchorsakLeftakTopakRight CaptionTemaTabOrder 
DesignSize�4  TLabelLabel7LeftTopWidthRHeightCaption   Gränssnitts&tema:FocusControl
ThemeCombo  	TComboBox
ThemeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder Items.Strings
AutomatiskLjus   Mörk     	TTabSheetPanelsSheetTagHelpType	htKeywordHelpKeywordui_pref_panelsCaptionPaneler
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPanelsCommonGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   AllmäntTabOrder 
DesignSize��   TLabelLabel1LeftTop� WidthTHeightCaptionVisa &filstorlek i:FocusControlFormatSizeBytesComboOnClickControlChange  TLabelLabel2LeftTop� Width`HeightCaption   &Inkrementell sökning:FocusControlPanelSearchComboOnClickControlChange  	TCheckBoxShowHiddenFilesCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight CaptionVi&sa dolda filer (CTRL+ALT+H)TabOrder OnClickControlChange  	TCheckBoxDefaultDirIsHomeCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption!   Standardkatalog är &hemkatalogenTabOrderOnClickControlChange  	TCheckBoxPreservePanelStateCheckLeftTopEWidtheHeightAnchorsakLeftakTopakRight Caption4   Kom i&håg panelens' tillstånd när session växlasTabOrderOnClickControlChange  	TCheckBoxRenameWholeNameCheckLeftTop]WidtheHeightAnchorsakLeftakTopakRight Caption&   Välj &hela namnet när filen döps omTabOrderOnClickControlChange  	TCheckBoxFullRowSelectCheckLeftTopuWidtheHeightAnchorsakLeftakTopakRight Caption   Välja med h&ela radenTabOrderOnClickControlChange  	TComboBoxFormatSizeBytesComboLeftTop� WidthlHeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.StringsByteKilobyteKort format   	TCheckBox!NaturalOrderNumericalSortingCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption0   Använd &numerisk sortering med naturlig ordningTabOrderOnClickControlChange  	TComboBoxPanelSearchComboLeft� Top� Width� HeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.Strings   Endast början av namnetAlla delar av namnetAlla kolumner    	TGroupBoxDoubleClickGroupLeftTop� Width�HeightJAnchorsakLeftakTopakRight CaptionDubbelklickTabOrder
DesignSize�J  TLabelDoubleClickActionLabelLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption'   &Operation att utföra vid dubbelklick:FocusControlDoubleClickActionCombo  	TCheckBox"CopyOnDoubleClickConfirmationCheckLeft Top-WidthTHeightAnchorsakLeftakTopakRight Caption,   &Bekräfta kopiera vid dubbelklicksoperationTabOrderOnClickControlChange  	TComboBoxDoubleClickActionComboLeftTopWidthlHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChangeControlChangeItems.Strings   ÖppnaKopieraRedigera    	TGroupBoxPanelFontGroupLeftTop<Width�HeightRAnchorsakLeftakRightakBottom CaptionPanel teckensnittTabOrder
DesignSize�R  TLabelPanelFontLabelLeft� TopWidth� Height4AnchorsakLeftakTopakRightakBottom AutoSizeCaptionPanelFontLabelColorclWindowParentColorShowAccelCharTransparentWordWrap	
OnDblClickPanelFontLabelDblClick  TButtonPanelFontButtonLeftTop,Width� HeightCaption   Välj tecke&nsnittTabOrderOnClickPanelFontButtonClick  	TCheckBoxPanelFontCheckLeftTopWidth� HeightCaption   Använd anpassad &teckensnittTabOrder OnClickControlChange    	TTabSheetCommanderSheetTagHelpType	htKeywordHelpKeywordui_pref_commanderCaption	Commander
ImageIndex
TabVisible
DesignSize��  TLabelLabel3LeftTopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaptionV   Inställningar på den här fliken gäller endast för Norton Commander-gränssnittet.ShowAccelCharWordWrap	  	TGroupBoxPanelsGroupLeftTop&Width�HeightcAnchorsakLeftakTopakRight CaptionPanelerTabOrder 
DesignSize�c  TLabelLabel8LeftTopWidthtHeightCaptionVal av &utforskarstil:FocusControlNortonLikeModeCombo  	TCheckBoxSwappedPanelsCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption6   B&yt paneler (lokal till höger, fjärr till vänster)TabOrderOnClickControlChange  	TComboBoxNortonLikeModeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeItems.StringsAldrigBara musMus och tangentbord   	TCheckBoxTreeOnLeftCheckLeftTopEWidtheHeightAnchorsakLeftakTopakRight Caption(   Visa &katalogträd vänster om fillistanTabOrderOnClickControlChange   	TGroupBoxCommanderMiscGroupLeftTop� Width�HeightMAnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�M  TLabelLabel10LeftTopWidth^HeightCaption&KortkommandonFocusControlExplorerKeyboardShortcutsCombo  	TCheckBoxUseLocationProfilesCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption7   &Använd platsprofiler istället för katalogbokmärkenTabOrderOnClickControlChange  	TComboBoxExplorerKeyboardShortcutsComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeItems.Strings	CommanderUtforskaren    	TGroupBoxCompareCriterionsGroupLeftTop� Width�HeightJAnchorsakLeftakTopakRight Caption   Jämför katalogkriteriumTabOrder
DesignSize�J  	TCheckBoxCompareByTimeCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   Jämför efter &tidTabOrder OnClickControlChange  	TCheckBoxCompareBySizeCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption   Jämför efter &storlekTabOrderOnClickControlChange    	TTabSheetExplorerSheetTagHelpType	htKeywordHelpKeywordui_pref_explorerCaptionUtforskaren
ImageIndex
TabVisible
DesignSize��  TLabelLabel4LeftTopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaptionM   Inställningar på den här fliken gäller endast för utforskargränssnittetShowAccelCharWordWrap	  	TGroupBox	GroupBox2LeftTop&Width�Height6AnchorsakLeftakTopakRight CaptionVisaTabOrder 
DesignSize�6  	TCheckBoxShowFullAddressCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption2   Vi&sa den fullständiga sökvägen i adressfältetTabOrder OnClickControlChange    	TTabSheetEditorSheetTagHelpType	htKeywordHelpKeywordui_pref_editorCaptionEditor
ImageIndex
TabVisible
DesignSize��  	TGroupBoxEditorPreferenceGroupLeftTopWidth�Height|AnchorsakLeftakTopakRightakBottom Caption   EditorinställningarTabOrder 
DesignSize�|  	TListViewEditorListView3LeftTopWidthdHeightAnchorsakLeftakTopakRightakBottom ColumnsCaptionEditorWidth�  CaptionMaskWidthF CaptionTextWidth-  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnDataEditorListView3Data
OnDblClickEditorListView3DblClick	OnEndDragListViewEndDrag
OnDragDropEditorListView3DragDrop
OnDragOverListViewDragOver	OnKeyDownEditorListView3KeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddEditorButtonLeftTop9WidthSHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddEditEditorButtonClick  TButtonEditEditorButtonLeftpTop9WidthSHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickAddEditEditorButtonClick  TButtonUpEditorButtonLeft"Top9WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownEditorButtonClick  TButtonDownEditorButtonLeft"TopXWidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownEditorButtonClick  TButtonRemoveEditorButtonLeftTopXWidthSHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveEditorButtonClick    	TTabSheetIntegrationSheetTag	HelpType	htKeywordHelpKeywordui_pref_integrationCaptionIntegrering
ImageIndex
TabVisible
DesignSize��  	TGroupBoxShellIconsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionWindowsskalTabOrder 
DesignSize��   TButtonDesktopIconButtonLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   Skapa en ikon på skrivbor&detTabOrder OnClickIconButtonClick  TButtonSendToHookButtonLeftTop8WidtheHeightAnchorsakLeftakTopakRight CaptionB   Skapa genväg för överföring i utforskarens '&Skicka till'-menyTabOrderOnClickIconButtonClick  TButtonRegisterAsUrlHandlersButtonLeftTopgWidtheHeightAnchorsakLeftakTopakRight Caption)   Registrera för att hantera &URL-adresserTabOrderOnClick RegisterAsUrlHandlersButtonClick  TButtonAddSearchPathButtonLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption7   Lägg till sökvägen till WinSCP i miljövaribeln PATHTabOrderOnClickAddSearchPathButtonClick  TStaticTextShellIconsText2Left+TopTWidthJHeightHint   För att lägga till genvägar, som direkt öppnar webbplats, använd ikonkommandon i 'Hantera'-menyn i dialogrutan inloggning.	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionAssociera ikoner med webbplatsTabOrderTabStop	    	TTabSheetCustomCommandsSheetTag
HelpType	htKeywordHelpKeywordui_pref_commandsCaption	Kommandon
ImageIndex	
TabVisible
DesignSize��  	TGroupBoxCustomCommandsGroupLeftTopWidth�Height|AnchorsakLeftakTopakRightakBottom CaptionEgna kommandonTabOrder 
DesignSize�|  	TListViewCustomCommandsViewLeftTopWidthdHeightAnchorsakLeftakTopakRightakBottom ColumnsCaptionBeskrivningWidthU CaptionKommandoWidth�  CaptionL/FWidth#  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowHint	TabOrder 	ViewStylevsReportOnDataCustomCommandsViewData
OnDblClickCustomCommandsViewDblClick	OnEndDragListViewEndDrag
OnDragDropCustomCommandsViewDragDrop
OnDragOverCustomCommandsViewDragOver	OnKeyDownCustomCommandsViewKeyDownOnMouseMoveCustomCommandsViewMouseMoveOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCommandButtonLeftTop9WidthbHeightAnchorsakLeftakBottom Caption   &Lägg till...StylebsSplitButtonTabOrderOnClickAddCommandButtonClickOnDropDownClickAddCommandButtonDropDownClick  TButtonRemoveCommandButtonLeftTopXWidthbHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveCommandButtonClick  TButtonUpCommandButtonLeft"Top9WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCommandButtonClick  TButtonDownCommandButtonLeft"TopXWidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCommandButtonClick  TButtonEditCommandButtonLeftTop9WidthbHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickEditCommandButtonClick  TButtonConfigureCommandButtonLeftTop9WidthbHeightAnchorsakLeftakBottom Caption&Konfigurera...TabOrderOnClickConfigureCommandButtonClick    	TTabSheetDragDropSheetTagHelpType	htKeywordHelpKeywordui_pref_dragdropCaption   Dra & släpp
ImageIndex

TabVisible
DesignSize��  	TGroupBoxDragDropDownloadsGroupLeftTopWidth�Height6AnchorsakLeftakTopakRight Caption   Dra && släpp nerladdningarTabOrder 
DesignSize�6  TLabelDDFakeFileEnabledLabelLeft#Top,WidthYHeight5AnchorsakLeftakTopakRight AutoSizeCaption�   Tillåt direkta nedladdningar till vanliga lokala mappar (t.ex. Window Explorer). Tillåt inte nedladdningar till andra destinationer (ZIP-arkiv, FTP, etc.). Använd Dra && släpp skaltillägg, när det är tillgängligt.WordWrap	OnClickDDLabelClick  TLabelDDFakeFileDisabledLabelLeft#Top� WidthZHeight6AnchorsakLeftakTopakRight AutoSizeCaption�   Möjliggör nerladdningar till valfri destination (vanliga kataloger, ZIP-arkiv, FTP, etc.). Filer laddas först ner till en temporär katalog och flyttas därefter till destinationen.WordWrap	OnClickDDLabelClick  TLabelDragExtStatusLabelLeft#Top`Width_HeightAnchorsakLeftakTopakRight CaptionDragExtStatusLabelShowAccelCharOnClickDDLabelClick  TLabelDDDrivesLabelLeft#ToptWidth� HeightAutoSizeCaption7   Tillåt att filer släpps till dessa &nätverksenheter:FocusControlDDDrivesMemo  TRadioButtonDDFakeFileEnabledButtonLeftTopWidthlHeightAnchorsakLeftakTopakRight Caption4   Bestäm mål för släpp genom att dra en &falsk filTabOrder OnClickControlChange  TRadioButtonDDFakeFileDisabledButtonLeftTop� WidthdHeightAnchorsakLeftakTopakRight Caption$   Ladda ner filer via tillfällig mappTabOrderOnClickControlChange  TPanelDDFakeFileDisabledPanelLeft"TopWidth;Height
BevelOuterbvNoneTabOrder
DesignSize;  	TCheckBoxDDWarnLackOfTempSpaceCheckLeft TopWidth;HeightAnchorsakLeftakTopakRight Caption)   &Varna vid otillräckligt med diskutrymmeTabOrder OnClickControlChange   TMemoDDDrivesMemoLeft"Top� WidthQHeight=Lines.StringsDDDrivesMemo 
ScrollBars
ssVerticalTabOrder    	TTabSheet
QueueSheetTagHelpType	htKeywordHelpKeywordui_pref_backgroundCaptionBakgrund
ImageIndex
TabVisible
DesignSize��  	TGroupBox
QueueGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Överföringar i bakgrundenTabOrder 
DesignSize��   TLabelLabel5LeftTopWidth� HeightCaption)   &Maximalt antal samtidiga överföringar:FocusControlQueueTransferLimitEdit  TLabelQueueKeepDoneItemsCheckLeftTop� Width� HeightCaption*   Visa avslutade överföringar i kön för:FocusControlQueueKeepDoneItemsForComboOnClickControlChange  TUpDownEditQueueTransferLimitEditLeft0TopWidthIHeight	AlignmenttaRightJustifyMaxValue       �@MinValue       ��?AnchorsakTopakRight 	MaxLengthTabOrder   	TCheckBoxQueueAutoPopupCheckLeftTop� WidthqHeightAnchorsakLeftakTopakRight CaptionC   Visa bakgrundsöverföringarnas prompt &automatiskt vid inaktivitetTabOrder  	TCheckBox
QueueCheckLeftTopJWidthqHeightAnchorsakLeftakTopakRight Caption$   &Överför som standard i bakgrundenTabOrder  	TCheckBoxQueueNoConfirmationCheckLeftTopzWidthqHeightAnchorsakLeftakTopakRight Caption1   I&ngen bekräftelser för bakgrundsöverföringarTabOrder  	TCheckBoxQueueParallelCheckLeftTopbWidthqHeightAnchorsakLeftakTopakRight Caption3   &Använd flera anslutningar för enkel överföringTabOrder  	TCheckBoxEnableQueueByDefaultCheckLeftTop2WidthqHeightAnchorsakLeftakTopakRight Caption$   &Aktivera köbehandling som standardTabOrder  	TComboBoxQueueKeepDoneItemsForComboLeftTop� WidthaHeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.StringsAldrig15 sekunder1 minut
15 minuter1 timmeAlltid    	TGroupBoxQueueViewGroupLeftTop� Width�HeightcAnchorsakLeftakTopakRight Caption   KölistaTabOrder
DesignSize�c  TRadioButtonQueueViewShowButtonLeftTopWidthqHeightAnchorsakLeftakTopakRight CaptionVi&saTabOrder   TRadioButtonQueueViewHideWhenEmptyButtonLeftTop-WidthqHeightAnchorsakLeftakTopakRight Caption   &Dölj ifall tomTabOrder  TRadioButtonQueueViewHideButtonLeftTopEWidthqHeightAnchorsakLeftakTopakRight Caption   &DöljTabOrder    	TTabSheetStorageSheetTagHelpType	htKeywordHelpKeywordui_pref_storageCaptionLagring
ImageIndex
TabVisible
DesignSize��  	TGroupBoxStorageGroupLeftTopWidth�Height`AnchorsakLeftakTopakRight Caption   Inställningar för lagringTabOrder 
DesignSize�`  
TPathLabelAutomaticIniFileStorageLabelLeft� Top.Width� HeightActiveTextColorclWindowTextIndentHorizontal IndentVertical InactiveTextColor
clGrayTextOnGetStatus%AutomaticIniFileStorageLabelGetStatusAlignalNoneAnchorsakLeftakTopakRight AutoSize  TRadioButtonRegistryStorageButtonLeftTopWidthhHeightAnchorsakLeftakTopakRight CaptionWindowsre&gistretTabOrder OnClickControlChange  TRadioButtonAutomaticIniFileStorageButtonLeftTop-Width� HeightAnchorsakLeftakTopakRight Caption&Automatisk INI-filTabOrderOnClickControlChange  TRadioButtonCustomIniFileStorageButtonLeftTopDWidth� HeightAnchorsakLeftakTopakRight CaptionA&npassad INI-filTabOrderOnClickCustomIniFileStorageButtonClick  TFilenameEditCustomIniFileStorageEditLeft� TopBWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialog#CustomIniFileStorageEditAfterDialog
DialogKinddkSave
DefaultExtiniFilter*INI-fil (*.ini)|*.ini|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist ClickKey@AnchorsakLeftakTopakRight TabOrderTextCustomIniFileStorageEditOnChangeControlChangeOnExitCustomIniFileStorageEditExit   	TGroupBoxTemporaryDirectoryGrouoLeftToppWidth�Height� AnchorsakLeftakTopakRight Caption   Temporär katalogTabOrder
DesignSize��   TLabelLabel6LeftTopWidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption?   Ange var nerladdade och redigerade filer ska sparas temporärt.ShowAccelCharWordWrap	  TRadioButton DDSystemTemporaryDirectoryButtonLeftTop-WidthhHeightAnchorsakLeftakTopakRight Caption%   &Använd systemets temporära katalogTabOrder OnClickControlChange  TRadioButton DDCustomTemporaryDirectoryButtonLeftTopEWidth� HeightCaption   Använd den här &katalogen:TabOrderOnClickControlChange  TDirectoryEditDDTemporaryDirectoryEditLeft� TopAWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogText2   Välj katalog för temporära dra && släpp filer.ClickKey@AnchorsakLeftakTopakRight TabOrderTextDDTemporaryDirectoryEditOnChangeControlChange  	TCheckBoxTemporaryDirectoryCleanupCheckLeftTop� WidthhHeightAnchorsakLeftakTopakRight Caption.   &Rensa gamla temporära kataloger vid uppstartTabOrderOnClickControlChange  	TCheckBox%ConfirmTemporaryDirectoryCleanupCheckLeft Top� WidthXHeightAnchorsakLeftakTopakRight Caption   &Fråga innan rensningTabOrderOnClickControlChange  	TCheckBox$TemporaryDirectoryAppendSessionCheckLeftTop^WidthhHeightAnchorsakLeftakTopakRight Caption3   Lägg till &sessionsnamn till temporära sökvägenTabOrderOnClickControlChange  	TCheckBox!TemporaryDirectoryAppendPathCheckLeftTopwWidthhHeightAnchorsakLeftakTopakRight Caption5   Lägg till f&järrsökväg till temporära sökvägenTabOrderOnClickControlChange  	TCheckBox$TemporaryDirectoryDeterministicCheckLeftTop� WidthhHeightAnchorsakLeftakTopakRight CaptionH   Behåll tillfälliga kopior av fjärrfiler i &deterministiska sökvägarTabOrderOnClickControlChange   	TGroupBoxOtherStorageGroupLeftTopVWidth�Height5AnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�5  TLabelRandomSeedFileLabelLeftTopWidthVHeightCaption   Sl&umptalsfröfil:FocusControlRandomSeedFileEdit  TFilenameEditRandomSeedFileEditLeft� TopWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogKinddkSave
DefaultExtrndFilter4   Slumptalsfröfiler (*.rnd|*.rnd|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för slumptalsfröClickKey@AnchorsakLeftakTopakRight TabOrder TextRandomSeedFileEditOnChangeControlChange    	TTabSheetTransferEnduranceSheetTagHelpType	htKeywordHelpKeywordui_pref_resumeCaptionTolerans
ImageIndex
TabVisible
DesignSize��  	TGroupBox	ResumeBoxLeftTopWidth�Height{AnchorsakLeftakTopakRight Caption@   Aktivera överföringspaus/överför till temporär filnamn förTabOrder  TLabelResumeThresholdUnitLabel2Left� TopGWidthHeightCaptionKBFocusControlResumeThresholdEdit  TRadioButtonResumeOnButtonLeftTopWidthIHeightCaptionA&lla filerTabOrder OnClickControlChange  TRadioButtonResumeSmartButtonLeftTop-Width� HeightCaption   Filer stö&rre än:TabOrderOnClickControlChange  TRadioButtonResumeOffButtonLeftTop]WidthIHeightCaptionA&vaktiveraTabOrderOnClickControlChange  TUpDownEditResumeThresholdEditLeft-TopCWidthTHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@TabOrderOnClickControlChange   	TGroupBoxSessionReopenGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption   Automatisk återanslutningTabOrder TLabelSessionReopenAutoLabelLeft"Top0WidthRHeightCaption   &Återanslut efter:FocusControlSessionReopenAutoEdit  TLabelSessionReopenAutoSecLabelLeftTop0Width'HeightCaptionsekunderFocusControlSessionReopenAutoEdit  TLabelSessionReopenTimeoutLabelLeftTop� WidthnHeightCaption   &Fortsätt återansluta i:FocusControlSessionReopenTimeoutEdit  TLabelSessionReopenTimeoutSecLabelLeftTop� Width'HeightCaptionsekunderFocusControlSessionReopenTimeoutEdit  TLabelSessionReopenAutoStallLabelLeft"Top� WidthRHeightCaption   Å&teranslut efter:FocusControlSessionReopenAutoStallEdit  TLabelSessionReopenAutoStallSecLabelLeftTop� Width'HeightCaptionsekunderFocusControlSessionReopenAutoStallEdit  TLabelSessionReopenAutoIdleLabelLeft"TopcWidthRHeightCaption   Å&teranslut efter:FocusControlSessionReopenAutoIdleEdit  TLabelSessionReopenAutoIdleSecLabelLeftTopcWidth'HeightCaptionsekunderFocusControlSessionReopenAutoIdleEdit  	TCheckBoxSessionReopenAutoCheckLeftTopWidthkHeightCaptionA   &Automatiskt återanslut session, om den bryts under överföringTabOrder OnClickControlChange  TUpDownEditSessionReopenAutoEditLeft� Top+WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder  	TCheckBoxSessionReopenAutoIdleCheckLeftTopHWidthkHeightCaption<   Automatiskt återanslut session, om den &bryts medan inaktivTabOrderOnClickControlChange  TUpDownEditSessionReopenTimeoutEditLeft� Top� WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@	MaxLengthTabOrder
OnGetValue SessionReopenTimeoutEditGetValue
OnSetValue SessionReopenTimeoutEditSetValue  	TCheckBoxSessionReopenAutoStallCheckLeftTopzWidthkHeightCaption0   Automatiskt återanslut session, om den &stannarTabOrderOnClickControlChange  TUpDownEditSessionReopenAutoStallEditLeft� Top� WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder  TUpDownEditSessionReopenAutoIdleEditLeft� Top^WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder    	TTabSheetUpdatesSheetTagHelpType	htKeywordHelpKeywordui_pref_updatesCaptionUppdateringar
ImageIndex
TabVisible
DesignSize��  	TGroupBoxUpdatesGroup2LeftTopWidth�Height}AnchorsakLeftakTopakRight CaptionAutomatiska uppdateringarTabOrder 
DesignSize�}  TLabelLabel12LeftTopFWidthsHeightCaptionAutomatisk kontroll&period:FocusControlUpdatesPeriodCombo  TLabelUpdatesAuthenticationEmailLabelLeftTopWidth� HeightCaption6   &E-postadress behörig för automatiska uppdateringar:FocusControlUpdatesAuthenticationEmailEdit  	TComboBoxUpdatesPeriodComboLeftTopCWidthbHeightStylecsDropDownListAnchorsakTopakRight TabOrderItems.StringsAldrigDagligVeckovis
   Månadsvis   	TCheckBoxUpdatesShowOnStartupLeftTopbWidthHeightAnchorsakLeftakTopakRight Caption-&Visa information om uppdatering vid uppstartTabOrderOnClickControlChange  TEditUpdatesAuthenticationEmailEditLeftTop&Width HeightAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeOnExit"UpdatesAuthenticationEmailEditExit  TStaticTextUpdatesLinkLeftTop*Width:HeightCaption   Läs merTabOrderTabStop	OnClickUpdatesLinkClick   	TGroupBoxUpdatesProxyGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption
AnslutningTabOrder
DesignSize��   TLabelUpdatesProxyHostLabelLeft"Top[WidthUHeightCaption   Proxy &värdnamn:FocusControlUpdatesProxyHostEdit  TLabelUpdatesProxyPortLabelLeftTop[Width?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlUpdatesProxyPortEdit  TUpDownEditUpdatesProxyPortEditLeftToplWidthbHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrder  TEditUpdatesProxyHostEditLeft"ToplWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextUpdatesProxyHostEdit  TRadioButtonUpdatesProxyCheckLeftTopEWidthmHeightAnchorsakLeftakTopakRight Caption   A&nvänd proxyserverTabOrderOnClickControlChange  TRadioButtonUpdatesDirectCheckLeftTopWidthmHeightAnchorsakLeftakTopakRight CaptionIngen &proxyTabOrder OnClickControlChange  TRadioButtonUpdatesAutoCheckLeftTop-WidthmHeightAnchorsakLeftakTopakRight Caption)   Detektera &automatisk proxyinställningarTabOrderOnClickControlChange   	TGroupBoxUpdatesOptionsGroupLeftTop� Width�HeightQAnchorsakLeftakTopakRight Caption
AlternativTabOrder
DesignSize�Q  TLabelUpdatesBetaVersionsLabelLeftTopWidthvHeightCaption+Kontrollera ifall det finns &betaversioner:FocusControlUpdatesBetaVersionsCombo  	TComboBoxUpdatesBetaVersionsComboLeftTopWidthbHeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TCheckBoxCollectUsageCheckLeftTop1WidthHeightAnchorsakLeftakTopakRight Caption"   Tillåt &anonym användarstatistikTabOrderOnClickControlChange  TButtonUsageViewButtonLeftTop-WidthbHeightAnchorsakTopakRight CaptionVisa &statistikTabOrderOnClickUsageViewButtonClick    	TTabSheetCopyParamListSheetTagHelpType	htKeywordHelpKeywordui_pref_transferCaption	   Överför
ImageIndex
TabVisible
DesignSize��  	TGroupBoxCopyParamListGroupLeftTopWidth�Height|AnchorsakLeftakTopakRightakBottom Caption   Överför förinställningarTabOrder 
DesignSize�|  TLabelCopyParamLabelLeftTop� WidthbHeight5AnchorsakLeftakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamLabelClick  	TListViewCopyParamListViewLeftTopWidthdHeight� AnchorsakLeftakTopakRightakBottom ColumnsCaption   Beskrivning förinställningarWidthd Caption
AutomatiskWidth(  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnCustomDrawItemCopyParamListViewCustomDrawItemOnDataCopyParamListViewData
OnDblClickCopyParamListViewDblClick	OnEndDragListViewEndDrag
OnDragDropCopyParamListViewDragDrop
OnDragOverCopyParamListViewDragOver	OnKeyDownCopyParamListViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCopyParamButtonLeftTopWidthSHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddCopyParamButtonClick  TButtonRemoveCopyParamButtonLeftTop?WidthSHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveCopyParamButtonClick  TButtonUpCopyParamButtonLeft!TopWidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCopyParamButtonClick  TButtonDownCopyParamButtonLeft!Top?WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCopyParamButtonClick  TButtonEditCopyParamButtonLeftpTopWidthSHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickEditCopyParamButtonClick  TButtonDuplicateCopyParamButtonLeftpTop?WidthSHeightAnchorsakLeftakBottom Caption&Dubblera...TabOrderOnClickDuplicateCopyParamButtonClick  	TCheckBoxCopyParamAutoSelectNoticeCheckLeftTop^WidthbHeightAnchorsakLeftakRightakBottom CaptionS   &Meddela när överföringsinställningarna automatiskt använder de förinställdaTabOrderOnClickControlChange    	TTabSheetWindowSheetTagHelpType	htKeywordHelpKeywordui_pref_windowCaption   Fönster
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPathInCaptionGroupLeftTop� Width�Height^AnchorsakLeftakTopakRight Caption   Sökväg i fönstertitelTabOrder
DesignSize�^  TRadioButtonPathInCaptionFullButtonLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption   Visa &lång sökvägTabOrder   TRadioButtonPathInCaptionShortButtonLeftTop,WidthiHeightAnchorsakLeftakTopakRight Caption   Visa &kort sökvägTabOrder  TRadioButtonPathInCaptionNoneButtonLeftTopCWidthiHeightAnchorsakLeftakTopakRight Caption
Visa &inteTabOrder   	TGroupBoxWindowMiscellaneousGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize��   	TCheckBoxMinimizeToTrayCheckLeftTopWidthiHeightAnchorsakLeftakTopakRight CaptionN   &Minimera huvudfönstret till aktivitetsfältets statusområde (systemfältet)TabOrder OnClickControlChange  	TCheckBox&ExternalSessionInExistingInstanceCheckLeftTop-WidthiHeightAnchorsakLeftakTopakRight Caption>   Öppna nya externa initierade sessioner i &befintliga fönsterTabOrderOnClickControlChange  	TCheckBoxKeepOpenWhenNoSessionCheckLeftTop]WidthiHeightAnchorsakLeftakTopakRight CaptionA   &Håll huvudfönstret öppet när den sista sessionen är stängdTabOrderOnClickControlChange  	TCheckBoxShowTipsCheckLeftTopuWidthiHeightAnchorsakLeftakTopakRight Caption&Visa tips vid uppstartTabOrderOnClickControlChange  	TCheckBoxShowLoginWhenNoSessionCheckLeftTopEWidthiHeightAnchorsakLeftakTopakRight CaptionO   &Visa inloggningsdialogrutan vid start och när den sista sessionen är stängdTabOrderOnClickControlChange   	TGroupBoxWorkspacesGroupLeftTopWidth�HeightuAnchorsakLeftakTopakRight Caption
ArbetsytorTabOrder 
DesignSize�u  TLabelAutoWorkspaceLabelLeft-Top-WidthzHeightCaption&Standardnamn arbetsyta:FocusControlAutoWorkspaceCombo  	TCheckBoxAutoSaveWorkspaceCheckLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption'Spara &automatiskt arbetsyta vid avslutTabOrder OnClickControlChange  	TComboBoxAutoWorkspaceComboLeft-Top=WidthLHeightAnchorsakLeftakTopakRight DropDownCountTabOrderOnClickControlChange  	TCheckBoxAutoSaveWorkspacePasswordsCheckLeft-TopWWidthLHeightAnchorsakLeftakTopakRight Caption#Save &passwords (not recommended) XTabOrderOnClickControlChange    	TTabSheetSecuritySheetTagHelpType	htKeywordHelpKeywordui_pref_securityCaption	   Säkerhet
ImageIndex
TabVisible
DesignSize��  	TGroupBoxMasterPasswordGroupLeftTopWidth�Height\AnchorsakLeftakTopakRight Caption   HuvudlösenordTabOrder 
DesignSize�\  TButtonSetMasterPasswordButtonLeftTop3WidtheHeightAnchorsakLeftakTopakRight Caption   Ä&ndra huvudlösenord...TabOrderOnClickSetMasterPasswordButtonClick  	TCheckBoxUseMasterPasswordCheckLeftTopWidthdHeightAnchorsakLeftakTopakRight Caption   An&vänd huvudlösenordTabOrder OnClickUseMasterPasswordCheckClick   	TGroupBoxPasswordGroupBoxLeftTopjWidth�Height4AnchorsakLeftakTopakRight Caption   SessionslösenordTabOrder
DesignSize�4  	TCheckBoxSessionRememberPasswordCheckLeftTopWidthdHeightAnchorsakLeftakTopakRight Caption1   Kom ihåg &lösenord under sessionens varaktighetTabOrder     	TTabSheetIntegrationAppSheetTagHelpType	htKeywordHelpKeywordui_pref_integration_appCaptionApplikationer
ImageIndex
TabVisible
DesignSize��  	TGroupBoxExternalAppsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionExterna applikationerTabOrder 
DesignSize��   TLabelPuttyPathLabelLeftTopWidth� HeightCaption    &PuTTY/Terminal klient sökväg:FocusControlPuttyPathEdit  TLabelPuttyRegistryStorageKeyLabelLeftTop� Width^HeightCaptionPuTTY registernyc&kelFocusControlPuttyRegistryStorageKeyEdit  THistoryComboBoxPuttyPathEditLeftTop&WidthHeightAnchorsakLeftakTopakRight TabOrder OnChangePuttyPathEditChangeOnExitPuttyPathEditExit  	TCheckBoxPuttyPasswordCheck2LeftTopSWidthaHeightAnchorsakLeftakTopakRight Caption?   &Kom ihåg sessionslösenord och överför det till PuTTY (SSH)TabOrder  	TCheckBoxAutoOpenInPuttyCheckLeftTop� WidthaHeightAnchorsakLeftakTopakRight Caption)   &Öppna automatiskt en ny session i PuTTYTabOrder  TButtonPuttyPathBrowseButtonLeft/Top$WidthKHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickPuttyPathBrowseButtonClick  	TCheckBoxTelnetForFtpInPuttyCheckLeftToplWidthaHeightAnchorsakLeftakTopakRight Caption2   Öppna &Telnetsessioner i PuTTY för FTP-sessionerTabOrder  TStaticTextPuttyPathHintTextLeft� Top=WidthqHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  THistoryComboBoxPuttyRegistryStorageKeyEditLeftTop� WidthjHeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrderOnChangeControlChange    	TTabSheetNetworkSheetTagHelpType	htKeywordHelpKeywordui_pref_networkCaption   Nätverk
ImageIndex
TabVisible
DesignSize��  	TGroupBoxExternalIpAddressGroupBox2LeftTopWidth�Height� AnchorsakLeftakTopakRight Caption*   Inkommande FTP-anslutningar (aktivt läge)TabOrder 
DesignSize��   TLabelLocalPortNumberRangeLabelLeft� TopxWidthHeightCaption      TRadioButtonRetrieveExternalIpAddressButtonLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption/   Hämta extern IP-adress från &operativsystemetTabOrder OnClickControlChange  TRadioButtonCustomExternalIpAddressButtonLeftTop-WidthiHeightAnchorsakLeftakTopakRight Caption%   Använd &följande externa IP-adress:TabOrderOnClickControlChange  TEditCustomExternalIpAddressEditLeft-TopCWidth� HeightTabOrderOnClickControlChange  	TCheckBoxLocalPortNumberCheckLeftTop^WidthiHeightAnchorsakLeftakTopakRight Caption    Begränsa lyssnings&portar till:TabOrderOnClickControlChange  TUpDownEditLocalPortNumberMinEditLeft-TopuWidthRHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       �	@Value       ��?AnchorsakTopakRight TabOrderOnChangeControlChangeOnExitLocalPortNumberMinEditExit  TUpDownEditLocalPortNumberMaxEditLeft� TopuWidthRHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       �	@Value       ��?AnchorsakTopakRight TabOrderOnChangeControlChangeOnExitLocalPortNumberMaxEditExit   	TGroupBoxConnectionsGroupLeftTop� Width�Height5AnchorsakLeftakTopakRight CaptionAnslutningarTabOrder
DesignSize�5  	TCheckBoxTryFtpWhenSshFailsCheckLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption-   När SFTP-anslutning av&visas, portknacka FTPTabOrder OnClickControlChange    	TTabSheetPanelRemoteSheetTagHelpType	htKeywordHelpKeywordui_pref_panels_remoteCaption   Fjärr
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPanelsRemoteDirectoryGroupLeftTopWidth�HeightcAnchorsakLeftakTopakRight Caption   FjärrpanelTabOrder 
DesignSize�c  TLabelRefreshRemoteDirectoryUnitLabelLeftPTopEWidthHeightCaptionsShowAccelChar  	TCheckBoxShowInaccesibleDirectoriesCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   Vis&a oåtkomliga katalogerTabOrder OnClickControlChange  	TCheckBoxAutoReadDirectoryAfterOpCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption:Uppdatera auto&matisk katalog efter operation (CTRL+ALT+R)TabOrderOnClickControlChange  	TCheckBoxRefreshRemotePanelCheckLeftTopEWidth
HeightAnchorsakLeftakTopakRight Caption   Uppdatera fjärrpanel varj&eTabOrderOnClickControlChange  TUpDownEditRefreshRemotePanelIntervalEditLeft TopCWidthKHeight	AlignmenttaRightJustify	Increment       �@MaxValue      <�@MinValue       �@	MaxLengthTabOrderOnChangeControlChange    	TTabSheetPanelLocalSheetTagHelpType	htKeywordHelpKeywordui_pref_panels_localCaptionLokal
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLocalPanelGroupLeftTopWidth�HeightcAnchorsakLeftakTopakRight CaptionLokal panelTabOrder 
DesignSize�c  	TCheckBoxPreserveLocalDirectoryCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption/   &Ändra inte tillstånd när du byter sessionerTabOrderOnClickControlChange  	TCheckBoxSystemContextMenuCheckLeftTopEWidtheHeightAnchorsakLeftakTopakRight Caption   Använd filsystemets snabbmenyTabOrderOnClickControlChange  	TCheckBoxDeleteToRecycleBinCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption!&Ta bort filer till papperskorgenTabOrder OnClickControlChange    	TTabSheetLanguagesSheetTagCaption   Språk
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLanguagesGroupLeftTopWidth�Height|AnchorsakLeftakTopakRightakBottom Caption   SpråkTabOrder 
DesignSize�|  TLabelLanguageChangeLabelLeftTop]Width� HeightAnchorsakLeftakBottom Caption-   Ändringar börjar gälla efter nästa start.ShowAccelChar  	TListViewLanguagesViewLeftTopWidthdHeight:AnchorsakLeftakTopakRightakBottom ColumnsAutoSize	  DoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReportOnCustomDrawItemLanguagesViewCustomDrawItemOnSelectItemListViewSelectItem  TButtonLanguagesGetMoreButtonLeftTopXWidthdHeightAnchorsakRightakBottom Caption   Hämta &fler...TabOrderOnClickLanguagesGetMoreButtonClick    	TTabSheetEditorInternalSheetTagHelpType	htKeywordHelpKeywordui_pref_editor_internalCaptionIntern editor
TabVisible
DesignSize��  	TGroupBoxInternalEditorGroupLeftTopWidth�Height� AnchorsakLeftakRightakBottom CaptionVisningTabOrder 
DesignSize��   TLabelLabel9LeftTop/WidthGHeightCaption&Tabulatorstorlek:FocusControlEditorTabSizeEdit  TLabelLabel11LeftTop_WidthUHeightCaptionStandard&kodning:FocusControlEditorEncodingCombo  	TCheckBoxEditorWordWrapCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Ko&rta av långa raderTabOrder OnClickControlChange  TUpDownEditEditorTabSizeEditLeftTop@Width� Height	AlignmenttaRightJustifyMaxValue       �@MinValue       ��?AnchorsakLeftakTopakRight 	MaxLengthTabOrderOnChangeControlChange  	TComboBoxEditorEncodingComboLeftToppWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight 	MaxLengthTabOrderOnChangeControlChange   	TGroupBox	FontGroupLeftTop� Width�HeightvAnchorsakLeftakRightakBottom CaptionFontTabOrder
DesignSize�v  TLabelEditorFontLabelLeft� TopWidth� HeightWAnchorsakTopakRight AutoSizeCaptionEditorFontLabelColorclWhiteParentColorShowAccelCharTransparent
OnDblClickEditorFontLabelDblClick  TButtonEditorFontButtonLeftTopWidth� HeightAnchorsakTopakRight Caption   &Välj font...TabOrder OnClickEditorFontButtonClick  TButtonEditorFontColorButtonLeftTop1Width� HeightAnchorsakTopakRight Caption
   &TextfärgTabOrderOnClickEditorFontColorButtonClick  TButtonEditorBackgroundColorButtonLeftTopPWidth� HeightAnchorsakTopakRight CaptionStandard&bakgrundTabOrderOnClick EditorBackgroundColorButtonClick    	TTabSheetFileColorsSheetTagHelpType	htKeywordHelpKeywordui_pref_file_colorsCaption
   Filfärger
ImageIndex
TabVisible
DesignSize��  	TGroupBoxFileColorsGroupLeftTopWidth�Height|AnchorsakLeftakTopakRightakBottom Caption
   FilfärgerTabOrder 
DesignSize�|  	TListViewFileColorsViewLeftTopWidthdHeightAnchorsakLeftakTopakRightakBottom Columns  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowColumnHeadersShowHintTabOrder 	ViewStylevsReportOnCustomDrawItemFileColorsViewCustomDrawItemOnDataFileColorsViewData
OnDblClickFileColorsViewDblClick	OnEndDragListViewEndDrag
OnDragDropFileColorsViewDragDrop
OnDragOverListViewDragOver	OnKeyDownFileColorsViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddFileColorButtonLeftTop9WidthSHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddEditFileColorButtonClick  TButtonRemoveFileColorButtonLeftTopXWidthSHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveFileColorButtonClick  TButtonUpFileColorButtonLeft"Top9WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownFileColorButtonClick  TButtonDownFileColorButtonLeft"TopXWidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownFileColorButtonClick  TButtonEditFileColorButtonLeftpTop9WidthSHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickAddEditFileColorButtonClick     TPanel	LeftPanelLeft Top Width� Height�AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� �  	TTreeViewNavigationTreeLeftTop	WidthtHeight�AnchorsakLeftakTopakRightakBottom DoubleBuffered	HideSelectionHotTrack	IndentParentDoubleBufferedReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChange
OnChangingNavigationTreeChangingOnCollapsingNavigationTreeCollapsingItems.NodeData
�     6          ��������           E n v i r o n m e n t X 2          ��������            
I n t e r f a c e X ,          ��������            W i n d o w X 2          ��������            
C o m m a n d e r X 0          ��������            	E x p l o r e r X 2          ��������            
L a n g u a g e s X ,          ��������           P a n e l s X 6          ��������            F i l e   c o l o r s X ,          ��������            R e m o t e X *          ��������            L o c a l X ,          ��������           E d i t o r X >          ��������            I n t e r n a l   e d i t o r X 0          ��������           	T r a n s f e r X 0          ��������            	D r a g D r o p X 4          ��������            B a c k g r o u n d X ,          ��������            R e s u m e X .          ��������            N e t w o r k X 0          ��������            	S e c u r i t y X .          ��������            L o g g i n g X 6       	   ��������           I n t e g r a t i o n X 8          ��������            A p p l i c a t i o n s X 0       
   ��������            	C o m m a n d s X .          ��������            S t o r a g e X .          ��������            U p d a t e s X     TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelComponentsPanelLeft Top�Width!Height2AlignalBottom
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder  
TPopupMenuRegisterAsUrlHandlerMenuLeft8Top� 	TMenuItemRegisterAsUrlHandlerItemCaption
RegistreraOnClickRegisterAsUrlHandlerItemClick  	TMenuItemMakeDefaultHandlerItemCaption   Gör WinSCP &standardprogram...OnClickMakeDefaultHandlerItemClick  	TMenuItem!UnregisterForDefaultProtocolsItemCaptionAvregistreraOnClick&UnregisterForDefaultProtocolsItemClick   
TPopupMenuAddCommandMenuLeft� Top� 	TMenuItemAddCustomCommandMenuItemCaption    Lägg till &anpassat kommando...OnClickAddCustomCommandMenuItemClick  	TMenuItemAddExtensionMenuItemCaption   Lägg till &utökning...OnClickAddExtensionMenuItemClick    TPF0TProgressFormProgressFormLeft�Top#HelpType	htKeywordHelpKeywordui_progressBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	OperationClientHeight#ClientWidthhColorclWindow
ParentFont	OldCreateOrder	PopupModepmAutoPositionpoOwnerFormCenterOnHideFormHideOnShowFormShow
DesignSizeh# PixelsPerInch`
TextHeight 	TPaintBoxAnimationPaintBoxLeftTopWidth Height   TPanel	MainPanelLeft2TopWidth.HeightDAnchorsakLeftakTopakRight 
BevelOuterbvNoneParentColor	TabOrder 
DesignSize.D  TLabel	PathLabelLeft TopWidthHeightCaptionFileX:ShowAccelChar  
TPathLabel	FileLabelLeft8TopWidth� HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelTargetLabelLeft TopWidth$HeightCaption   Mål:ShowAccelChar  
TPathLabelTargetPathLabelLeft8TopWidth� HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TProgressBarOperationProgressLeft Top*Width.HeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder    TPanelTransferPanelLeft2TopKWidthBHeight?AnchorsakLeftakTopakRight 
BevelOuterbvNoneParentColor	TabOrder
DesignSizeB?  TLabelStartTimeLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00ShowAccelChar  TLabelTimeLeftLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00ShowAccelChar  TLabelTimeLeftLabelLabelLeft TopWidth-HeightCaption	Tid kvar:ShowAccelChar  TLabelCPSLabelLeft� TopWidthAHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption0 KB/sShowAccelChar  TLabelTimeElapsedLabelLeft� TopWidthAHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption00:00:00ShowAccelChar  TLabelBytesTransferredLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption0 KBShowAccelChar  TLabelLabel3Left� TopWidthBHeightAnchorsakTopakRight Caption   Förfluten tid:ShowAccelChar  TLabelStartTimeLabelLabelLeft TopWidth3HeightCaption
Start tid:ShowAccelChar  TLabelLabel4Left TopWidthYHeightCaption   Bytes överförda:ShowAccelChar  TLabelLabel12Left� TopWidth"HeightAnchorsakTopakRight Caption
Hastighet:ShowAccelChar  TProgressBarFileProgressLeft Top%Width.HeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder    TPanelToolbarPanelLeft2Top� Width.HeightAnchorsakLeftakBottom 
BevelOuterbvNoneParentColor	TabOrder TTBXDockDockLeft Top Width.Height	AllowDragColorclWindow TTBXToolbarToolbarLeft Top DockModedmCannotFloatOrChangeDocksDragHandleStyledhNoneImages	ImageListParentShowHintProcessShortCuts	ShowHint	TabOrder ColorclWindow TTBXItem
CancelItemCaption&CancelX
ImageIndex ShortCutOnClickCancelItemClick  TTBXItemSkipItemCaption   &Hoppa över den här filen
ImageIndex	OnClickSkipItemClick  TTBXItemMinimizeItemCaption	&Minimera
ImageIndexShortCutM�  OnClickMinimizeItemClick  TTBXItemMoveToQueueItemCaption   Fortsätt i &bakgrunden
ImageIndexShortCutB�  OnClickMoveToQueueItemClick  TTBXSubmenuItemCycleOnceDoneItemCaption   När operationen är klarDropdownCombo	Hint3   Åtgärd som ska utföras när operationen är klar
ImageIndexShortCutF�  OnClickCycleOnceDoneItemClick TTBXItemIdleOnceDoneItemCaption   &Förbli inaktivChecked	
ImageIndex	RadioItem	OnClickOnceDoneItemClick  TTBXItemDisconnectOnceDoneItemCaption   &Koppla ifrån session
ImageIndex	RadioItem	OnClickOnceDoneItemClick  TTBXItemSuspendOnceDoneItemCaption   &Försätt datorn i viloläge
ImageIndex	RadioItem	OnClickOnceDoneItemClick  TTBXItemShutDownOnceDoneItemCaption   &Stäng av datorn
ImageIndex	RadioItem	OnClickOnceDoneItemClick   TTBXComboBoxItemSpeedComboBoxItem	EditWidthnHint   Hastighetsbegränsning (kB/s)
ImageIndexShortCutS�  OnAcceptTextSpeedComboBoxItemAcceptTextOnClickSpeedComboBoxItemClick	ShowImage	OnAdjustImageIndex!SpeedComboBoxItemAdjustImageIndexOnItemClickSpeedComboBoxItemItemClick     TPanelComponentsPanelLeft Top� WidthhHeightnAlignalBottom
BevelEdgesbeTop 	BevelKindbkFlat
BevelOuterbvNoneTabOrder  TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeft(Top�   TPngImageList	ImageList	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
u  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ��JA���.��v�R��E!�+d/��
�]hu�+T��EY7]iu�T�P bAY�nQ�;әugYM��\,;3��۝���9tSD !p�iDe���d�� �+�1��]���D�4˶W<u= �C����+c'%�\���Y;R����
���)�(K�eHU"3�b;n" Ҽ��@q\�,(6�+,I@&�дx!�5�k���ƪ�!Dӵ�aJ���-
E�Ͻ1v�7�x��b���k�!B�a4`P �#�󶙟��r��( �$���:p��h�p���L��6@�� Ҭ�y
��i��ၸ �6kh��� �}�t [��f}���㔺�g���CV p-�am?U�m��OI�h^P�Ź�*��c�#Äw��$�(���?(�v̢U���!��2�z��eB�)��8X3פY��T|Z�0�Ŀ��\�n�mB���,    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   %IDATx�c���?%�qԀQ�����xM�g��t �47� OWL    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
@  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڅ�kHSa��������nnS�v��0��D�҇>d����.�>!+��KE�A*]i؇AHV�(���9�S�e��gz֙et:b�/�����>��%�eY�����?m�}�%�F�>Ռ��,V"���7�YK��U�E�29�$&gcO�N�q��}���b@�eJ�^�k+�L1?G��@G� &���s��+!lN�Z���g�,$󽴝6`�������w$��C�U�yV���h�RB�
�n��� Oo7�a$q���R�]pzb�|��$I�~��B9�514���8|qk#�6(�z
եj��Bj1�����?��Ds`)1���oA�k-q�xĄ!^_���q�}O�����,�G�C ���6r~�qȍ9𴖒17պ<��u���Y"/�UT6|D��������R�H4�>_��.b>� lw��YݥPj�i�
�r����Y�4.���͋���Ez��-F�F�#I(Y��f@�(�f��Q���aD�h,��W���L%�YUC�8���'���2�m�������\+����߾�0���DZb6	_���U��E�AYo�ji�_�����V�A����L�|�f�Y2	�d
���É_S���-�Ҟ��A���_�|�	v�J�?�����^��    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
g  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڍ�[H�qǿu���ߦn��.��l���H��z�2H�6����zﭢ���$�A�`�0H"��4��x7�s�9us��o��T�����9_>�|��f�mKTr9u������b���:���<�s/3��N�(E�$� O@G�^�����W��������v@�3�镤���e�1ŜT\�FV���}����*��2_��8]�/��zy� C����[�87Ϻ��lkUS�N�3�g(rKI>(Rpq_+���.;��4�[����<�������<#��P����.�0,��]��*z 3��RJIT���{�Pood��@m�%*� �Mc; X�4e�F-�ݚL���5�@�1)�u.�M�=*��<�"�v��ko$y�C�$�
	��F�'nO�3?��=�ж�&J]������O>���:����_)ar1�A[!õ�����N���p�`&�#��1��ؽfM��|)��V������y||����` ��^\�ЇKr���Čs�	��g)��G�z��+b�KdF.��qa�)_}_?�Kq>�{h���mi��p���e��3O��1a..��^��z�seW���Wf(C���7���x$	UCvǈͶV�+��H8^������y��$!1qMO|��r������HRE%rZ�!������=(ZD�0L�_Y�'���    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
o  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڅ�mHSQ��ws���n�l��tS�Hi(�2� ��T؋Zm�!�L�}�@VЇ�Do�I��K�/���'M�(�R��t�D�:���IB7��p��9�w��<�!���͡z��� `�V��X��,���)�c�)��A'!;d�Ȕp���\[YƂgޥ��L�wt����v@�fRԣ�6�Fhbx��(db��c��q~q��#!�r�"��6n/�����\�j7\?�aui��D}�S�>��Ů�ۗFJ�<�1N��fZ��xd[�ڪ����;�
�� s�rl�Q.x��j�&�p�z?���c��/��b��z5�"S�w�#����F<�s~\����������֧�hp�l��~�q��:f��5���#6(��gFY�M3K�;V���V��q�JK�
yQ�d�����A�4���B�P�Ķv8�����f�n��r.a8��dcú劈T�\	s�W�h��»J+�>�"�d���)P��������{z��`��F�����TB�O3(i4���A��|]]���c�f���!��4� �#	�,�8��ʕm�á�0x�0e< ��B�V�=�WE��O�E��h�H���}�}}��~�B����x~;�Z!����33�ij�@���wq콽p��]\�H-E}�
��U�q�n��(�V�o �����'��~��[w�h    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
2  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڍ�mHSa��w5��ۜ�6��K�
D���L2���|k#��^�/�)
�(*��ERD(аr�A�L
�	BE9tw+3��ܜ�n��g�I7���{9�=���s�s
1�`L��R,d����w��v�G��+8�y�:3�-����)���ʨs~��{�ٙ�|0��u�zb1 �gZ:�N7�j3E��4)��lc��d��@���L(��z�IJ��3��I-�k&5XZ�����Y�QGGy�(�h�e��ӌB�1$�Y�͇���}��ƶ�o�V�>;G!�HD��]���co�n<��e���E�̕�F���d��� ��x�i�[]������8 R�:ݘ_���ŚL�Oq���C�4���^�v>FxjT`&�g�p����s8�����)���:X�Ԩ+M��C$�ҳo൑�yY�Q�@�
�� �ۿ�p~��+�L�7iA�<�HJ�c*����߮�á�8����B�N�������θ����Q4HRZ�+c�`d4���UP�g��(Eg�.j���'�T�Ʉ׫j%���FY�l5,AJ�E�>j�y�v�B�P���Q��_�ӆ�e��x4����K���k\`2���	�1��S�W�����_�$��d�E��?��'������    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
U  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥSkH�Q=����cM�h����_|?�F�@�R�勘3!C+�Vj�Y*LK,4QDJ41��&�A�E�{d����oKMt�r/�q��sϏ�&�d��d�R bP߳I���R��蟝R���>��
����=AA�G򲩴�$DF�{δZ�g����sb2�{ͺE�J����z<���z�����i��/�e5��w�v8�E0ň��;���q�^����C�*��ޛ�VYw�$8�;@�ALN��Nz��=�F�QЈ���|5����H��)�����n�>�]�V��|>��|8�	�~�O�~�w�O417
FI$�:���E@��r�O/�)���4�%�]�P\R����u��&0��@4j��eP�7��A���Qu^o$�<ä�!�w1;;���8TV�##=�K�v�����˨����+����s�he�B|f���r,,| �����l6�Y�� �-�ɕ((<m\#���lX��h������"22m-׼:�������{	V%�D?��3V\'`u	�db��X!4�ZW%xM,:��c����,]k�k���y m"�B#�8�?���|c(�;/�J�0��Ό�)���
�=�pON��3����dEgl�9i)�`�o �oh��is��U��>`�Xp����(�j���d��������� �QN�^#a�    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  PIDATxڕ�]H�Q���5g6�B�}�]A��$e�[�Zi�MW}X�Y�UX�E$�^�F�J��E��L��̹i&��bm��u��w/��6X��������A�Sq��Ʈ��_nn��Z�Gx���c�/���q"7��w�^��/@H"�ke�P!ߊd�3C�)�����q�$��/���9����dL���!�^��D]?��eY�2��˄�gdt�]���@�d)�7�F{��Lmm��.���o�=1\k���QSg )���2�p^��O�.��D���[X�7�Jt�Q�	RvSO�+���B��L��c3B4 ��z���Q�pRK�X��'@NiZ)�,�E�+j��H-@�')SaO����$�c���@N^J�*��``��ڵ&�0�L�*
c�?���	�~瀔����꣨l��9�g�n�>�p $���q��"mz;����\m���NOt�m��0��_ D@V� 8wۮtU
�P��Q��8�M����q�?�u{� ǪS��?c$ة�AqH��!�>/L���u����)R6�Y[��Z�h,F���a��W�Z� l�OFCL�    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  DIDATxڕ�[H�a����G̠(���r5�Eu�%!���,o���C&�i�	l��[�e�hjih�eЪ!�d����m���>(���ދ�9������ZM��}�`$�Q�7���B��WZi��D���a�z��v�Bѽ<�,F5cu:Jr�I��9�b�냽cd,�M��|=�K�{���a* -��>������n�?~z<�'@��j��&mv�֡��ȩ'�U�l,1���TJ����Q}����Cj6�⌹��pm�.��bA�2p�]5����5�h&ȉ:e� ��ox����$��vF�����AՐ�����'��洁�h��)��
~������a�a+Tr$b���cn�c�-��8��p<%�ߵ��(|�^��� ?�C�=}Rt�>�T���*%@�хn�dB)W�&� �A�/�A���G��|�g�4߀�uk�VA!S�̉��5!��f}���VݥL�a�����u�t#}����ṁ3;�U�ը�(��%�͜�BL�p�#�G�\�U�`����F�)`�k�뗟��D�䛬)O�w�H�ɸ�[�����#�� �    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��o�d  �IDATx�u�KLQ�l�bR|��<�4�D�Eqa��2F�5��hD�RڢF4j\��Ђ�%%���A6 jx�h�<RJ��ӡe:�X�C���{n���s.u�a;AРz���A��z���6��xa�����a����^��"ԅ{�H퍓py|����°ɂ�O���re�ifE����+?�ku�+Պ�� ��f8�����٩"���Ud�uyEi�L-��c�W�P"���f�S�⺮�"cO,�;�Ѡ�%7���4l�8T�#N����Z�B7��P?m�su�W#�@" _)Euѫ�Q��
 ��lD����X@���%�P��/5�K@|M$Y��U�yM�U�:�+H�o�>�~�Ʀ��6a�,�j*@X�z��<�3U�D�.��a����$˓"��G|��,��X���Z��5Ld|8�LP��D�.��	 Gc'�	%	�y�6���e|�E%�@�2�
�D�Q`Ʊd6�bK�L�7��>ɲ/,&m3��Y@�׋��@�;vo�����{�^�JC���0�M@���H~M�i;A�����8="���J{ǿG�{$�]C�)ObȮ��v�;�j�<��6-����gu ���Q���x\1��&�����?H�wz�:E-�^��    IEND�B`�  Left(Top� Bitmap
      TPngImageListImageList120HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڭ�[K�@�l�]�-H+��"���`�C�L�'��"�~�}�/�"�eETD�n����&�g�,�$��K6�s~�ٙ94�"�
�RښXw�/�g������l�������mɹ���NaѢ�r��0��U��Ұ�Ba�0�����piޫ�$@����#����Jl������  �m�����5�g�Y��ކaU��h����Z���Jm�	n�����O5PGŽ�=��|�[�Vn�,�>��p��;뙬"�(C��$"�y��~kIT�Of��V u�;�Ģ��*:
�KC� ;J�^� ���� ��Jl8g�%�z�_.Y`��!`�
V�E�;J�Eb�%�CbY$bd>ӷ���6v	mJ����2N �;���nlq�,�"�n��5�_i%�*z���8.@|��=���G�o4L]4�~ �p,Л�ھL��/�B�h�g�/9D��������3cղ�r���6���q�� �    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   -IDATx�c���?5㨁��8j�����H�@���5��^t �C�����    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
'  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  ~IDATxڍ�]lSe��oOK�Ӟ�]�֞J{�BƖ��8I\a�!����M���No�FB4c!Q.����$��1�Q�F�4���@YR��tY{66ۭ_��9�=�m��IN���s~����������K�쁢4��%(����H 8Acdlb�����t݄���n�����hu(�Ȧ�E6�~��Q荎�G6>����l�Y5��X�aiqn�����<�q�;o4�-6{Uб��F~X���������=��'���^������U��V-���I�{������8B6�<,��MT��?�R�8KU���-��\�������Z��,�$|oT�pqGK_@�!!��63���Wq%�R�K��f�4Cg5`��ӫ}��e�%E�_ia�ŀق�7?�+<o��� ���!/���Őώ�v3N����l��;���;I��$=��T*"&�J��[�J �aC���0�6����h��ȥ�h����q/�E�HH��c�\G�YV���ҙ�����pBT�.��>���5���{z���V���V��?� 9���at��ċ��Mf��)<��/],�}���_T
~�mβ�k4���w���,���$��CϾW���X1���W���WӹL�]m��l�M��f3������yL݉C"g t΢�ujY���Bg�M���EwQ���69���h �2���ZX��	�d2���[�c��v�C/�*�.z��ڏ�{�%e]nfW�L˛G<1a�*���u���1�ܾ�lx���������\3F�K綘�E ����匕�Kf�����;�,�{�z�h5�V'U`#�^�B���J��TZ)�}�P��*��z�'t8����,(�2��<*�X�/����RG�J�,    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڕ�mlSU����]�{�vݺ�ŮK3��	c��h�D4j�L��$�([H�~ A�ň�@Ld�ė����"1dq,s��$V�vs�ۺ��-w�����V�8_�s�s��<��s�;Fi��<��fdd����	���*{r�� n�-=v����h���2+�l1(��$e ����MA���E�ԑ���o���mN���r���C�L^�"����=�d�w��Z��`�(zc#K1�=�'�����G�w���|���ϣ�qGmU�
¬F_�i�Ǟ�a$�&�^���_t�.z�~P�n�q����7���atb;}�|.��U��r"�s?W��ɇ����,Y$}�K��8N�����$b���)�B[!�h�v�74E@���x�S��Z* �2^�Ăx۲�G𹉂Z+�Ec��O�f��~���^�%�}r���÷~�f%���p���e)P��lۤ�rxg����
�=�Cح�)��� �@䲐Ij�!��M���,knO����{l�Z��1�W���m��q%{[Z<��������sb"���cA�4|���tqܮ�rSg,<ݑ����<g(sit���V�ᮟ�S_�EKO+^tِ�S�f�?m:�3���������X�����:^�s�*qz��H��m{Ƃ�\?��"%d��\�gQ�X���1��?#@�V9�8��/��fO��R������c�Z]W����� I�\bf��ƑC����j��Hj��ՠ��7?3۰H��vE~��W�٬\�zeѢ�!e��Á��=�߷�a2Y *�;�D�f�O�x�����*�<��b�cUhE��،H$^�Ƨ�z `�FcW���-5Uk(
��3sI�ו4�%�	a����}�~���+f���sJ������JH��G8�a,}M�d���_!��|�fv��rRX�>ߞN�Z�²k$���)�d~{0���rcm���� M�/�����"���\��    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڍ�kLSg���=�^�U�)m	�Ʉd�lj&�Z��f6��\25q�b��1�d���/[�h@�b Ǿ�Yb���)C-��,��9�={{61�bx�����������Rx"��,n����l+Dq=(jb�H�ܘ��N���L�V�d�U���u&��k ���|3��H<�y��9�V7�T����z�Z㊷�NE0��x��;+ ���ݥ�rM�-:�!#����q�-�`z2���׃�߷f�O�7t8U��ٶ)#̔C�7r���($R��F">�7���}9���C��԰���׫t����Z�;����|l�d�Wo��ؕ)�p^A�)݀e�����k�8�=�|��|R�'�3yK��~4A�)IQ?W��g�$x�?b�\��]�1C�u�I.���0��b->h���8>�3J�}s8�]:�L
�����r ��3��*5��kM�Q�M2Z:#h&�i9�t6�X�X�����
���H�(��p���BPZ�]
��U��A�{�ނm���Ms����!/�{��0��(��5�1#�Ja4��'�)GS<���C��~�խ��4��B��,b%���(ں�p���� ��$~�	y�A�6�@�B��]�
B<��RQ��:�b�l�^�$��Цj#��.̠���2t	��=�=��^'����{e�0���������Ĉ �Y�R���F��EZ�(S�X0Y
Ȉ��Tnvp�(��WL66���[�1V�	��ۑ��G�SY�+<7�����������,�7r��5C5CS��=-yO��l�q���e>�g���J&�Rx�*�����Қ����GV�p ���Y�~��rAG�5u�mp~?�X�ŗ�%���w�쪀��J+��n�i����w�)*?4��-���u�e��KV���K�\�n��5i��;O��9$]o�������J����e�&Hw�a^�y�������� \�&��    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
B  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڝ�mL[e��OoKi�-e��ގҎ,�e��e!˜����e��\���/�$j���t�[�����[�\
���[��vMB����е�������:�e!���<��s��=+��䰶�@d� �� d�0*|�s��h���w�Z]&E��O�����9�5�`�
��)$bQDn�X���I�%���{ ��/��Z��!ê_����T��͜�Ϭ<"�qԍVp��:}UAг�XJ�f��A���:�V�|R��ߢ*a{��G
¸29�>W!�[>	a1!`v�w$�wx�����i��%�� ��.�X���x�9/�b����A�Ӿ�P��յ[�� �^�ޗ��k��:�o�1ɟI��O��y�F���C��3�t~�V��۫��E�{ϋe�~���n�8�`��y�0rt٫��f��	�GO�${h�.��re2i��Ќs�!H{���جR�x�iM�Z�!pl �./g���^��% &#�W�	O �E��bvu�Ӽx���^	hr\hU*�.}�z��S�&4l��/-�B�� .LB���X��o���b�N�_���T���>62����f���+��J�C;���0+�/��Ű��G���|�\	>>�Z�H�'<���O�d2�Yj���~�X�1V���ҳ����R� 6�2?��WM���J�9�l�-�Lv�T�pY��� W*�U,EJ�d2� ��!]dd�瞒tV�%8^��g������B��c�/T�}�W��H�g�(�)s���CB^P!����;n��l��ޚ���k�����r��wg\��k�o�c�+��4Xڧ�r�O6���kGG�(�eM@)�Ǜ� �K�iNvٰqC)�sK�|=�st���ֱ���5�bݹۢ$�7 q��T��^���1�>`i�-�P    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  +IDATxڍ�PTU��wqw�?Fa��݀0h�����V�lR1����U�aQ�&,²����r���Z���P�V�0wY����{(
�y�9w���y��-fIX�CDH H8��^
b`o=8Է���m�#�|G��WY`Y�R�::�9����.���2t?]�=���v뛿m�?�(,*�L敝�s;BW-���o C}�c#��T���A��9��+?��p�P[˹<��2X�R��ٓ���ZA-V`�6�����ӠA*��WC{�=��<4g�62n���w�Ѣ�p�� r�*(��(�A��A�@G���y�
9L�2���Æ[	m��o��T�}
>X��u4׈ ?Wx:�bzM8/�#BXu�t�6~�
j�����V�`o����H£�_cRk�5�_�cF��~FpX$�޶>>��6�8�}����ri*�����}j��?��w6ǭ�����I��q�fh166����Hھ+W�υv�
�V�1y1�(?~�K>���KV�u ��i),��DҎdLLL��bT((ȇ�Tz_=�z˒x-�!���9�����J'K�{���|1�/Ĵw\®�t�l3�[R|P ?0�Ph{+ ��z��o�yO ֜�r򠵀�!����٠�8���pvr���SX�l�C�v8�Ex�����'d ӣ��fI�r�3� �!�H:�dۖ��������)iق�3i)ɛ� ��X�L.����a1�-`���w���B�:����&8HQ[�I���ڙb{X\7�U�0�l�T�K�ɍ� �kD~u~��J;<ڱ��P�*Dvvw�`s
��=b���U�+�H����D�>��xM.\>K6jK���25�[Ǹ�:L�b��)䇄Z�k��zX!���G����tmq)?J�pȜ3m�����W���n�R<�(���OT|rCC�#,3~�p󁂱1�&"r84$heĺp���&썎�	�_Z����5�9��M_?O:]�TJ<Wld�)!�
�U�	�����x�lOO������hFV��    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڝ�YLQ��k�@n���D�/>�
!��e��E�.��(��T�J4q�D�A(!�75"FA6�*�E�RZB���8�"�-��0wNν_�/��������)i���|yV����Yx�^���	̚r���s �u_��Y+tI��w����p�F��lZOC��@Ż�vп��B�Й�2n������t�aLk�7��M�B��������!\8W:�ch��Ε}�(L�"v��(�����	2w<h�FԾoEQj4!������D!�}��	OjP�. ĩb��p��j��=I���r�d�YL��MSY��*z�)޺>�7)�/�b�˫bد�xi��R}|�����=HyX�ҜXB�ߖ3��(�h�]Bg���e�6�`T7��cr<�5�,WLȹ��L�Y=�������rߖ�H!Lz f��y�b����Ĩʍ'�lN9#K`�29�z�.�<��a��I�V<�ʬ���ްX�ЫiPJ|��"�~��	�T��!�Z�����lU�>0{��۲f�	F�c�I�����I>9�Y���E��'���!� �34��/`�<l���Ƨ����LFOb�Ki�)�;O�?r&`bA���~v�C=���&�`�mb�Jiz,�NK�!4��<�[��}��f4[9��g��"I1�P�	��!0�p="�"�٠����/�t��*�6i(L.rr#۪�;��_	m)9hKs;:*n@�)Z��U@��'���Sf�}�Q�h�9��#��u؍�    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڝ�kH�Q��g�:/�%I3�2��>ERQ�'�K)�p^��]�Ke�獲$�O�:���kIby)1����;�ni��lSO�&ڜ�xy��9���w�C`�.eVR��Ǵ�O�"P�F�RK����iv�	h�su���H�>7O�4z蚀��4': j��ܔR��~9Jj�Z����I*L��)r\;{}�Ԉ��q�M���B��|���� -)����q_�X3h��;ٰ~��wyqA��Ei]�x<��ۏ�uC���O��-ݸrT�N��C҃r��	YU��U�2��_���Bt��I!�XR��i$u������kc�$x�J��;O){;��۰�E�����낃��_���pBΥK�8.��y��K�>�����;r��.$��*�স�J��Sڊ��uط� l�6`8�1���YY9���	9������sf�,Ш(�:�Oά-��0 #RѼD!b������w��ϝ^��tЪ�J�Tr1�B0�4�PWQ�RL�-S�c�nX��\]�� �ܤ0$�Ox���	հ�o��=�bt�����c�^���04���¡X%aTvzVp��f�q�a�u�0>:�����δ��� �/`F@>�5K��
���ߑ`��+�ߛff���l��8:�2T*��r�06��l���t��pv��Z��Q=L.5tj��2�3P�_l�����͆k�����Ym���t�i����^�    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
Q  �PNG

   IHDR         ��   	pHYs  �  ��o�d  IDATxڍ�kHSa���Q�b8EPԔ���
4�H32"/hZ��X^��!�NS�.� /V���H`i�i^�:��nz�sy������p������y��Əv��fIt}V��n�|t=D�5���N``l��-�ᄃ~����%-��d�:�覌� ���M*3#A3� �n0bR��_K����<{H�U�E���!���fCEj�)�}��a0��1����Q� �]�Ajn����v�l޴�J�:�_��.'F�Q�Jjs."���VyJ$��:ѐ+f<|Gjs/au���x�=	k��g$�s=�Q+mlGc�e�O"�7=N�^*M�H� ���
l[O��qx�Eqx�^���V4߉�G�ݠ5FP�-DZxJ=c�>񄟯/��e9��G�,�EKI�������\��H��_�fv2���/'o(i�il�@�Yp<�?cTU��Mp���2=�Ĳ���n���	#�����=��,a��]�bQ���,�,+Վ�A��T�P	�ψ�8����.>���p9[�i��B��V�7�#E��<]!_u���HK� �X'�y���9�lΥ^��rJ�q�=Cܰ0�_�D�JSl����9�as��*+����r
�}Nx`nH��A�"����q��
t���&,e�D=d�Cs�d�'~��B���
�'9��KL���t���Fz��OF˰���R����V���a�`���g�j{_xT>u���)��9�Oߞʲϵ�j�� �k� Mȝ�    IEND�B`�  Left� Top� Bitmap
      TPngImageListImageList144HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڽ��/�@�gZ�Ŷ��AB�F��"qw�pę�
w���_��]D"$B���b���ߩVf�3��Ի�����g��}Cc$Ϡ�&����U��#��2��ݗ��@���:%t�0���y5��ኂN���i:u����y��p���6�J�o|��Y.Ivl;��mk#>�G����>�z�K�_G�E׭5	�%k�l�sc(�#M"������_jx�`���A%��jY��Zb2!��Y5|!�M�W���p ݽ��+�Q2i�	9w��M�LA,)A2!I���S��� SKlHH�~��3�]�kܒ`\#8����-JVFpQr	��Hk��Ë��H� ��sW��H��״��1~��{$JAR n# �ΪQ����� �2h�ƻ  o���B: ���|��Rc�M�s�Gûb���ԋ����G$�]<�!pJh��\��G��!P�k�����@�#.J
���'�#3��]�#����    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   /IDATx���  �@�_�XȖV@�$�2� ��x~^��N�S�{���    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  ZIDATxڕ�kL[e����;��B[F)8��1.��N��bչ�AL�4�M4�~��b��s�xul]��l�m���D� �`�Ph����z=��D��u<''=�}�>����PH kw[�Q4��PNqM &@Q^h��҉�j�K�Nk!͡E*WlSg�@���I�{�H��\���u�챷[������
�e~^c(�j�r�a����NLO���hl��OϜO	0V)b)�E�y�V�R'UVHhH9���y�tG�������_c���5UhHX�����.ir���bx:����h��ղ5)�Tm��I�g�E���\�?�ľ���nw�w$H���#����Y�&����˫Ug��Z��q������D���\S���=�jy)�5ǯ�JJ$YR�k39|�W����tµ��\�Z�^�؃j�/��TE�tR@}U&v<�~��l3�=��a���m��%��-6*�V085���$CS������Ugu��+�����L5֡5��ui��4�7�[�K^4�¦uJ|�k!<��:����"��Ǉ��J*N�d��ZU���8�
����"D���@�1੏���-Ğ�� wA��q��r��b�&ۻޞe����8�$}_��-/@�fW�����8���OAi~�%�0��T(�`�9���~���!w���hjmv�\�����+f�.z"ʾol��^�gP{�e��,{[H��(�z���t~>��]�����^Mf��[,�i�3à��l{#� ������n|	��䩓���W;��E����)T�5���7T8���}�P�a&�	��f�������頯>R,��/��,�� zC3�B9�b�f�ƣO��L�q�t�#����u�I�a�%	�����[WXYUA%��E י��Ԛ�$�Ì��+�KeҔ��`���X�1㨩��\�>+��s�+�c���Q&Qr�7�In��.>�c��"�,x�=��P�j(�%���'���w�}A��UHwJLm+c�h�*�52������=Ax~D��[��:���(y���E5�!T&~ڈ�5���� 4��������d��8�j    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥVklSe~�9=�ڞ�-�z�ڭl$&b���`)���8'[%^�&��b"&j�ˆ��d��x	bw$���&�]ح�lmמ�[�~=����__����|����Ca��Y�ZN�T��(���%�PԩD<Qӵ�Y�\�?X\94�J�\�\�ˀ��B���\42����ޫ��#(�q��0@����i	�M�ٮ���ԔH$��_������Vu}���X��:$��9;_���)+�4d,��c(�Go�%_41:�]�p�ulŮ�z�m��<K��2�����il�b m��Ȥ�j籎*�Ҕ �"�RV&?bq���k�Jl^1��/��G�s�DFC�:��G��*v}�3XK�����Ā��8�m��X<!��}����Y�||j��L��3�Ҵ��3u,>/7�{W]��N��ᑤ�:�V�O͠��:�p4M�شB�u�U��ъt\O���8�[��j'���={`^�j���%���,h����Q��{R�$����H��n��e�@�y	\�g#9����>,�Ubۆ��y�{���O*!�q�5�N�K)2��SiI�����VL&A�l�hX�F��ؤ�8�}�E�*�/����F�0��O�aPK&<��+{��~��=p\:�ڕ��!��6���j��d�U�6r�ی�Y3��OX�Pk�/�+U� RTl̆q�Irm��gZ��u�+�n���aÏ�=�9��3�J��f���3rl�&�Ǐ�9��U�l�FgT���A@��fì���k�;�D�ٵ�f�����ũ�M��o.C������\�J�Մg�#~Axp�ٱ�w�S�)81&�2�@���	&��f���E,�3CC@z=���r:��=/{�%]�ӿ5%����f�;����I)�#F��-�sH��f�c1D�P���Zϕ�|Ͳ��eЫyty�!!�Z~i��>�`y� T�"O��uþ�hF����$�x��?�E����СJ�<�b%�YgHҘ�z���Bn�u��p��=���d��s��t�|L�&¤����, <�� ��������iˢ���L��hr��{hxky@�rK ��+iv��Z�F޽s8��A����(�\���Ax�#ϖ�޹i�J�s��sf9��p��бޠ����F���"e�O����pb -�i�U��i��2����G��c�����73������Ϸ�A���%6@m,���R�=C�s�+��X���֪�    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڕV}Lw~�zw�Уł���!�d�7>��͹�M�L��D�������c&�1�h��tS�P5:t����f0��R�@�*�
����Nd��7���}�>����9
�X��MeAS( B�@(�(�em�dVc�F=��e��Y�*U�K5�p�!`X��axh �v��#��86��e6� ���T�Q���5����}AE8�����2 x}�ڎ�{�"���2��ZDlbH�Z��p GC����t����c����<x&�)�\j0��%e�\I㧼P�*�?���g\f�gk�d9���/�)ۼ�U�j"�. ��ja�2���̎��QR.��܀�1w��Xf� sr�?��Q��Y�g6�4W��,#V��Oe������[�f~<=��SMƘ���<Z��H�Q�7�;Q|�>�xF�^ܱ}'qz�fg��j���f���`�~݁Xz=�1A�����z,��;`Q\ 4�
\ltɒT��[�@���.��OI X��@twvd\<K*�g`�i�na�n$�a��G��}���S���6�#J��ɤ�����q�n�A������&��x}���߇k�'��l�H�qa74�'R��)R��+.r��@e:Y�a��Г䥟�@�a�|ɟ�C��Ue�R�oU��P ��V���zI�,>F �؆\�v�
��',.kB�RUA� |�Ɋ~����N$�䩍�xI��:=������V" )����n��_�mr��*h�^�3h�	����y�����6����rY�T�#5  Ɗ
0�9qT��'& �d?�	�ח���.ћ2uٱ�Y5���e��S���
�s��o��r	���ٲ�iKd�c ")kk�����|3n���S��1�|G���X�RCbC�:�r$�]w<+�N�T����*C��"����^��M�Fh�m��9Ѩ�x:�]?QkO.��{��is��uq,CE74���k�;�Ի*�}Y9��ţ�f{�~{�Jyuǫg��kk�ص�3�͛�)*�]����^]1�a�O\���ۉ���45Mƹ�x.\��0���h�zO>�>^��S���C��#P-]����46�KHO��X`}c��:�Tь��.	��/�,���P�|�`�08��Sf����r�'
��<7�R	�.VQԆX�0�4�dy��	�'2}H����.��3r��� ����+(q��I&�1���[��|"������ܿ/*􊆗�!    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
   �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  wIDATxڕ�{L[Uǿ�����QXy��x�B�,�E^b��&���$�f�H�?�Y�C�0Q�L�9�tNp.�@4�<�T@�ĹQ��Q��M�z�-C:Z'iz�����߳��`�~I�B�T&8.�x@Q��U}�ր'��EP�.�fP*��SJ��{A�H�=�yK�x83����֌Õi�'�>V�@�E7}B�<�U䱔��anjFC�,k����[�̮�SҶ��h/����a����f�X,-�a��ެ�[;0R�ѻ- $G��
�x�8U.��e�7�e4
����h,�l(K;���;�He�FĂ��qx�+
Smֽ^9���U�.`D���J�@yZ�C@p��s�_P�b�߶�*��C���e�%c��� 83���/�Ҏ;� ��ou�޽��S廕��Ts]�����3�V�X�({!ڱٺ���X7���
R�H?�!�s/00i��cYý]���i�N�a1��r(�"�ܽ(�����;OW�y�N��q �o`������sa�K���<ީ��3{\�^��=�Q�6g��L
�8��O2)�i�I���<�H�Ӹ~:�����Cxk��b��>��U���a5�;GJ����7���7�������M��gI;h�Q�?����P�)�v/��{�+Fx�`�߁��TM r3#���bjf�w'QQӇ�����u�y
�O�hQx�$�\=�!\z5�uK�Qxu <X �w��o�ב۹��>�qn�X�����O:��
�k4��T)��t�'���0xI�5������[�S�����!9^m�;���j�}�c��ܕ
�� �IDBA�,��Po���-�@�+�^H�����OC�p��®;����$�H�$JenୡE"[:Z�`��@Y�J���|�k��
��ju�~��n<O��GH@�y�x�g�J8�-�譃��޵����s��v�m�x*Ik nP;�ۑN������j9�}���A]�0>(�#��I�8����o�ه��,:~�ƕ��F{�|�����s�F��t�:x����L~��T�ڎ111�2���f�HIT#?+
>JLN�
�|]����r�������ӎ��~�6�$0��`�kc �ۤS�t6ն<:�/����0��    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  nIDATxڕ�{PTUǿg���X\`�QAK�0B@(z���A�2��N1ڐ�H"�a�/�	
2���ZHj�-�q45ЕF���>�ν +�:3w��s��~��w~�A�_�Lw�D:�R�A�M@�)%v��@�$ '-sau��Gi���	�+���rAS�1���NN��&�u����
�5|[�� ����@} ��å�<gN��a�a`�f�$Δ�����ۑ_X����z�lz���T񀀀P�'G宄�d��8A
�o ��@�o���F3�������T�Bp��=lMI���u�e%{� ��5������-�u�$mZp7N �ZP�%l0��F�kvt[	xx��|�� ������� ����ّ������6�7@;;���l&] }�uM�X$@T0�ݽ�؄$���4����^����E�[�tQ4��u�<��i� �PP��4X<|@흻�nmn^ʋ@[�ۘ�R�5ɀ����%��B�j�;�MGG�����9��=��r����?T��Љ_[g��cP�8��} B�>$6���\��olhK�ׯ}-t���u��u܇�A�����ឋP(�`>FGA�T��4ԃ�a�!����O 2ve�|�/����ؘ�~�7����&`�aV����[���:vvv�1K��^Z�z2�ˊ��!Y�1*�^�����wg�s�n�m�1�D�ad4,��8t��e~�#&�˱�/1���J��~�*��D5���B���?��%���ּ�L��[�Y�ō���@�T|GZ:����S�g���	V�� ~�,P��2p�g��i@���ǲ�;��������철�aȻ\��Q�'�8�����Ϸ���WB���v���#6v�
�YϺ�� �"��������y/^���+&M�����sK6�d�H��[]��Ï�6�#`ʋ��+ �o	�37.C|j�����"�����HJI;�;L�ǰi+72��0L^�6�8����wE���e}2���/��tV)j�� �A�4�����O�S��&
�����Y;`V��@�;,і�C�Zuc�K����ya˗��Jr;l�r�<0���E��o�g�,�8�29y��/:Xu�dEO��:��n�,;�w��o;$���(�/v����ʩ0m{qQ9�?����؄7�'��ȫe���^�?X�R9����n8CB�ٖ�A�4��*/�x�ާe2K"e6���,ły�bl	%���z�����������6}��^%��mQ(����@��G�������X��ŕʫ�|�����#&cg�����W�_�����z��pH��u���Y�h��=����<)��T��@��y� u�s    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
S  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڵ�{Lw ��2P��+�.��ǜ�Ɍ`��q ���թ����h�!�[����h�hb�D#�t>��Z���*(����{��w'�;���e��������~��5�!�?J(��x���R���Y�V�V�����~[��p�O���כ_ɐ�.�B�O��h�Hk����^�z���/G�6�;�������ͅ�vכ^�ߥ�|�����6�ö�*a�n\kj�� �G/�`ϺYT�@4�<}�FA�d�b x!�����`-J�������Ɨ�8V:�E�FIu��3�@��������o�:�����T�"��зBx�Rm*���߸ �+/�r���T���_�(��	Y��؁2�IԔ.E��d��T��^PW��\���]u�ÙB$MH���͘t5$�PY^X�����~6�ݜ"pؾ��ʝ�JVIg�$M��!��:�螊������f�ib)�@q�9E�7C��cDW
��j��D�����
����؄A�~p�xq�����:	��<I,�s��b�i������o7#s|>4��.�7y�b��������>�_D�-Fg����8�mȁ�zV��/��Y��4�j����7S�F�и�3�=OX��.�5;�1LF��Y++�%�����(ɕ����"1L ^��	q=�!�C{��5&�������&k�!�͋a��*u�2��I�	be�R5 ]<����>�Q�)�e�
S�x�W��??f�������t���P.�K[�Rl��R��?#kn�,4��n���f��9���p�� ���A+� ��X�de+V���?w�U��&�AX�i���a+�sh,e/�`{������ 2 ����;?W��`U"r�����\����Վ�+�d�s�Z�0vZ����'�9�Ј    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  XIDATxڵ�kHSa��g��.��� �� �(Bꛮ̂.fEEf̨��B�T�Pt3�Y^"�(�\s�Q���Y3S�45ӲU�y����9��M�%��������{��y8�!��E���<nRfW��U5L�Ȭ�f�
��Upqo��].z��M�]$-�X���ڃ��F�U���9�¿����i("C0I$�������=&T7~j��b�G�/�T5v�ج8�tߏ�]��ӈ̃�(�_"���1e�6���4��{ϡNX���<��H��|��Js�r���r���[$��x�$-6̱?=[�줨�_"ig�1+�GB��ۗ��@z�y)�y���r)^�a�ͭ��D�mF~y;�Z��i+ذ�$h��P^}<�^{$���Պ%KC�'B � `����,�����h�Eq�C�e�ʡ�0[=6�v~��k<��*q쿬#���H̪�zrvJ�O��;"�(�_R��/�U�z����g�T�y=�:��`�R	�T�J�Z-/�s��h���T?�
��.Br�K,Y
Y@ #�����g�M�|�x�W7�zÀ���!�ɜ��%z��(N�%�c[qDU�n4:).��8��	>h����㙔=,��'
H��0L|��F#NެCPp��K׬�l��kC-�Ŕ��W��yALZ>Ѥ�D�J;����¬�� �Me�p�f�lBS}-hڲ��#������q9/؞r�h�w�i�䕾������H(rH~���`�X�э�7q��_d%}}�t{A�'�v4���n#b+W׌�W��oy�������vf��@��2�&�S30}f>��[�W�8�s����\�1E��1��XOp��l�:�pX    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
A  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  �IDATxڍ�{PUǿk�Q�@J�2@1�XV�NQ��T��E��^251.X�8	#ro��A�������:V#$�{�%��޽Ͻ�{Z��	�k������>��=�*<�3������d}^��.w���,i|�e9���ӏ��zauȆP���4}�
��u\�1�q������AS����ggHs�z�B��i���q��'�.�z���p��A��}�{7�Cx�� 	bd�uu���xcZP���v���Mpy��+��`B�u8~�;����U*(����DS���ﮄ~b<�� �ۋ���}[�v�N�e[��yY�g�q�P��Ek�����?n#��m�]�/�*^�u���u��j{p@�����"V'��0嘀@,^��'�a�i��	ȯ�R��"�9�ch��K�xD�i���0�ٙR�����;� �jc.�͚iM@z�<�)�U���O5�!"*�Ӌ��4T<W��E+�\iݷ8Q�{7��G�I�ð�vU� ��\��^4|��h��"9)�����"���P�D*�;p�<��E�v�ܠv��M�.��W��Y�����\�g���`�2!^����,�ٯ�D-Y i۸Ԏ�#��*Fqf�:} �$-K@�"�N���a�<���q)�Z���{�)�,zTNY+9��ǔ�/�*�����F���	�m�y�
7����n}��g�r��1ZAe�jIsUA@��G��_� ����s���ʀ��r�g����)7�o��DC�� ^:�c�#P� w�at�x=dmX8�W���^�� H\�.C��8�9�i��Z�\d��mz�V/���n#�_8�Җg<8w���tr�z�&D�c�����_��$�^�<���w�i���1³|�1����n��ϤJ��_���<�����M=̓���s��T�����%}��O���1p��g�`-5��| ��YOK���� ���#^������B�k�/R�2��x�]�1�����/M    IEND�B`�  Left� Top� Bitmap
      TPngImageListImageList192Height Width 	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
p  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���AkA����d���J����A�b+�ă'Q<�$��C꿰�
�Q�^s�x.��VDPPJբb�M6U�3��mv²�ٝ�:��fw�'�Lv��������@).��	%�R�����A&^.�/½"I�k�u���]�4@4��\ղ�z�]!��"0nS�lڶK���m!� b�������l;���"T|⣌���U�w������yW�q�q.}��j��k���������M`����������*9��5K���B�0��$���j=7��=/��.�b���� ��/�Ec��L�^�a����@TR&n�����5����5��(�փ �����DoA��[O��gm;�60�:vŇ�S�(� Zù�	����#�d 0��A�w�Ѐ{�s��N�� � x��>�E�
 ��[�e������g ��I��r�j�0�b ��OB���D����HAT��߀���'a]��L � � ~�#)������{��z�k?BD�\ <���1ƴ�O��q��q�"�ei���9lO@�f�q<���6�/�v+��#� j[B<��@R�d~�z|Ab��&�DM ���#:��Hԑsc�7N�O"�q ����{q�#Y�P:| }7�'����(�dr(M;��o���B������z�������F~ŏ    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   8IDATx���  1޿�	�Hz����Y           F�\Q�W � �����o��pf    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�ŖLSWǿ�����E�>h��F!�|��W\|L�(�	d.:�,!�fY�s�t1Y6c�e1s�tf>P�.�L&*���),��m�@)X
}�{{wn�l���&߹�|���w�w��1��0 ðI_*��V	9��وaLz�p)`�y�Cv��q�X���B4oT�h������b�,���< ��H?�]p9� E�=�e�������Y�JΦ �/��s���b�tf}�{�����qy�b۹B���.&384Hdqq�L�p8}������>�����[�}��=m 6�L� ���V� �(�1X�*��nl�44�[���y�+�E�H.�p��&����?�,�%�p�(��N_ E����&C���K/*����!I�a�T2���2�.��
�(
��]�xh��47b 4��8?�;�H�v�J�$A��JB�Ik�MQ(
��`�O��G�RR}U�Z�Ԇ'F���PJ����+v��kx\��#����#PݎR.U$�0O'��%��M���t�����?`��A�y�a��� J�]�tB%
p�@	+�G��5�����	}��6��wכ*���-Ai�]�I���M#@̓+���F�!�@͞�`
��c聆v�� ���:�A�<R��B�I<]���(�ؙ���^4�<� l\$��֏�~v��=�Ɋ�=:���A_@I�4xat\|����ّ��d���S]�5z6W+>;u�	T\�����{<�k���Y����)D��Θ�9j'�_������4-�kTP�jL�c��i*A�]x���A��,�|��2S�@�ւ�YN���^<�h�c�6@�e���� ����"!�U*W�	�,4H�Z5l{mb1�E�݊����6�C���	s2�#|�C�A���h��`����'�� ��I�Ue<.��\�\.�?�5�=?n��Wu��v�9��K��Z���A���B]}��d�ܮ�Cmc��A��x�/8����cKt�Z/Um�	[�lA���Aq9�,�AFjzD������7޻a�k_6��l7H�����Ic�(����)m^���;�k:� �Z�bʰO%v9���N���	�ֳbB���q��(B�nB�I��S��-0CjJʴU�����A��)�Uz�8Gлl�!��1�[�}�!oU2���8�N��y��s/��޺���2��~�BM
��.l�7����ݰ�M�p���ΰ SIw4f8��l n�ޞ9@�ј��K^�$DQ3p�<p�vӣ�D�{]F�;�D�}Y�v������, d+�Q���1�4���V��+g0!��MW��Ƈ�G��@�,m������Y$������F��C0?�8� �虣xfJ:"���pY�+��D�-FCV،�����l�9,���x'pϗ(	��	��IO����}n ��-?E���?�2��B F��y���)@A@W1L�t��h��Vչ���g}�x�L��"�    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�ŗlS��������G�W^$���A��QP˦J�B�P2:Z����Q	ZU��]�Ic�P׎D{tk<T
4�Q�mt��.�����ډ�'ر���^��\�z��(fDڑ,�s�w��;����;�$I���Q2 EQ~�?}���5k)�~���r2U@pEH�#+/��Q�g��������iҩ̶�%�ڡRk��
%yQH"���1%��%���/��N�3@i�{.@u�(������'],��a�߇tJ<�ǅ���Z�(��R&1hcMV�sFh��i!�@��*Q�-9|����ѻ��Θ�m�9������g�q�W@ �B:�Bwg;�D젷ٽ�����èt?+����N�j�Kf��'$�5�%���D:->��;�3�sS�]#Q]3�z�e�E��bώ7�v ��
r��qq�����9��?Ǩ���O�K{v�	�b3���~K�"��%ґx���	�U���1��h��hjb�w��nTd��Nq����>߿�r��=�=9Z���\��z�<%@u�����Hn���������C=���}����lj�ųuj�~J�]��X9gD��U��'�=�kv/���Z��f�(�f��4+q�RIq�^��4��,�\A������+:!��P����H� �-��
�Tk��\q���'�n"�L�����#�/G����1Q1#�'i:��y���Է$�k�ւ���on.�
�wǰ�?~C��/�d����m4�L�魛_�z��m��uN �u�?�dT��E��MYؾʁK�]	�r����}]�%�m(�$3 py�u{s��2�5�N����Lُ�W;����Ũ�X�����̩�aT^nE{�<�)t��5׬�H�n�v��KD��?��ɦ�uG�
���(�B��/Īl\n��Ϗ�q�B0;�ć��e\�!��4�T�]s��['&P�,`�߳������p�ϣ��n�����R=&����}u!�V�2�@X�S��N�r$�2�(ִl�|]T��+����A-K"��Q�UD�a�Ÿf���"8��qL9���1)�G
��6�ى%�Y�ˍ����{I�y����ފ�`��������#��m �`P�����Z�pb�>��"����=Hl��3��̟(�Z�ձ�%�NZS)�H�>�%�/cٷ�BŌ��ھ���[��%D��j��Ӗ7��Jē�^�@4�ص��^��MX����6���?�oĴ��/
	RxY������mݪը6/�w�j5����c0��8���rIh)|�~���^�ނ��r+�A�J���$�B	�H�~���q�墳�l#��ը�/.��V�!J�g�6���H�s�n �ǚ�"�gIL�s�����_T+���\%��u�9Y��.���I���(������%�sr~�C]l6f�H�������k[��+��`?˺�V;mL�A�	� �xqO��ӛ�H�S/4��7���~3C����Q6�H�����Qe1�� �	�g�<a�y>�7O��w�ػ���,_CҺ�(:y�[Jc'��Ag�Ib"H �	�v7��'���`X�������DW��AA���]~�`�"O�S.���B�A������Zy� MZ�(��S1�R�	����I���#ۢѶ1r��t�BQ>W�B/��H
�iqA�^/���{�����R���V���O��cYRդ�6����D�Ҵ��_�J�};��H]`P�X�y� �9*�%�    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  "IDATx�ŗ{LTWǿ�3�0/�d ŕ�	Fj�n����X[��֖>\Mt�]7٭�f�mvY�ݭЦ���Y�*�H�J+զ6T��"�2���0ܹw��s/ʊ"L�����9����9��8#�y�O� �d�Aӳ��*��X"�>-��S�++�e���h6�~�������?+�mi�Za0���%�J�F�O�J��LNd>�D0�#�	6�t�?:�^���M ��:P#�1�2��'=PY����F�'�([dJ�W������Р�''[&eC*���&B���z ���<�>V>��m����!)ǒ>�q����J4�xQp\�M`�����%�2����vJ��S��GcZ�[�$`�d%B4��J/�4GvbP��8v�ӱ�D� ��GL*^�f�4E�KWɬ�c�+����x�KvA�>O��W��.�3 Y�zJ����X��B=��֊�V��ݞ�(˒]�L:����%���QVsJ�d^�hJ���^������;O�P{)0bN����m���1�@M	��x�a\��tv���>K�~YE'��#ÿ�Ӊ@��3�㙕���	YR'��q����܄�9C��6���g=�͹�����>��[R����m��] yYjXr��@��j��[�b
��э���Q�}7ζ;J��
В`L�V�>�GR�P�>U�7uC.�#����K��_��������Փ4�s8%e��� �W�����j���IMal�Ӆ�w�RT�=_�D�Y;`�vI���A�҄�E��x%� ���
9�8hJ����)3V?�8<��C#ˬ~^��]}�����xݟ1�u)$�%�GQ�X�a��qp��:�Ly9M�� 0�:��W)Zu	F�Z�6�q���_���y��G�ov_Fщ7�(;�t�b��a;CK���Cn KJ����D�>b��<8? ����C�rU�`N�L&��SV�)L��P�_�A��²��1+�57�O>���8�{{Ź��dPYY��}���nAGu5.����#y���wU�m���ܣ�B�X���K��E6��1�}�-+��B�2�ŵ��<�def�z�sH��}�v�5@�b�wU�w	�uh���U��/�Q��8t:I|���ru�&��a��):�{��:w��{���&�V*a;[*'�＃�����wbؼ��[���q���َ �ϻ�Bb\Y�Q+�O%R��8��܄��Vǹ������EQ��A������ �����ܪ�D������~��0}͡�Qo��!��`�>(���Ol��A/&��]h_|=e�8yrL ��0�����f=��#��1/���>w$O.��Jm<x���t��"�T�r�0Ts��5s�c�<-����A�Ղ:�	�� ��i��(�ͱqO>	�c�`�����!�·���h�O@�m)PP�i۶C�a�6mB`��1u�ϭA�{�!�ԄV��\���S�u�3f����ׯ�=w���Fi\l�_A����;p�����N8���h�k������z�"�O����ep��H���0V}���%�Е�K���p+�=4��.h�M��gۍFXI��,�� �{7��Fq�r�thI���i��eh�p�,{�$��	�K��L)�͔��?�d+���7�@���^ōK����I*�yO*~8!�0���&��SIQ��A]\E6�ZR������8��H�Ѩ��\r_1��|�UN���H+���d�(���c�K�$���� ǝ#�^z-@����Y �Ȯ���B
'�#���n�p_���P�Խ:�B�?.�l��    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�Ŗ{L�W���7�}񒇨񱉈�l>pjE	N ӹ���d�\b2E]�?���IgDE@���M�?�(W��mAZ(�}~��WFgmi+��$M�������s1� ����0��h�Y1��Z�a��F�@C!�
t#���]M���(on3�Q����، ���3�,�/ �T �[-f�ð��6K72�RU�\P�O 2�|4 �-<W\~��Ƥ퀶�/T�۬��FK��B�a� QY�Q�\�@ �6(�O��MХT�i� 7�{�u�䍼6 �v:_$�ϑD�̋!��AR]�� �m�nk�i�\Y&�zm���K����ط|������˄a�'5`0��F;�[תd�>Hr+E,k�6����j$����OE�~։�"/����I��ceن�>���3�N���E>L�Cn
��n�@^q�c�f�"/4��@yV��'�蜪��`�{A�0������j��렺i�I�[�FGj�����jG)���
ɂ���mEY��H������C��*��;�VK�c�L?� 2D�bΘ�M�0���3�ӀN�ը*���v�U:ahL �%���l�Р�y�ֱz�fR�zw�=I�-�y��[ }ߋ�J�t�� ��°���`n����[�F��s5�>����~2�G���b�v��i�L%����SU����D��ض�R�z��t�Q46;�e;s���k�>���� ,��@1��L�p=G�{Ǌ���7��p�}i�θ 
��ea�j1d-r(���`����g�Cg���&�}��]�MYb`�|�~�9M�(�m�B�o���0���x޽?�ڝ D�8�,F/P(as��Ev����%���!��'EO�T�(E)1j�/M�@~�<�gӝlȓ��S�e�uf�uݽ��F ��Ӳ+�hT��@qP��� V���T���Wt�/�t h�D�q�����#I��2\�������:Ө%��ϫ�T(��q��F:/��]kB!;M8��Al��%�z�:�B����Z'�o�-r;WU��cŏn�o_Y�T����x<���N����'h��<Pj��30v����c����.��qlϿj��r��p�y�I/�(X���^B\��{V���#��y����D�s�J8Q�(��M��B
�+47e�?�A�d��Z
TˀG ��zh4��:��=>JI	��2�F%�ўg�n(��w	�%�1��EʋV@p �e�h�Az�5�W��$ai���x�;wr9�Xo`QZz+z�͜�|�YÓ�{ -�Gd�ݓ���A���$�s��(�x�� �&�i�WP1�O:{�!%q�4Tv�3i ���7 �ws�R��
O?j�{�6uJ ��+c)�Y;=�<]����\o1'�rON��J��Ԛq��"ػ�m�r\�Q�u5-Q�-&�Z�b4IX�jF���s�[�1�A$`��^��Z�P����j�����q�7�8��U+�j�,��!Ծs����ᶊ����������qA`�    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  mIDATx��WP����,���]Lg��`��7h2iY�4
�0Z3h�P|���HŌ�cD�Tl�;�Heq&�G	�|�j�����{���Jw0�ə���ݹ���s�e8�Ï)�a�q,]$T�����爪�a�'vZ��
,W^�6��,R�c��0�C*a��J��ys���4L�Q��Ã�����w�h�q5u��66����YZmŃ�0_��r�,���j%|��
k{G'N���T���W����D���a�q�۾3Ȏi��`�4 -W��@�=p&�&<����#�	]�D"�y0������[�_�� `�T�'��k��J���I`�}`�] n\������l� ��,��sT��(`�������F�x�F]�8� ��I�7���B� l�l�	��ș�Ѱ��}���"0�w3�Ltv��๑K@l@�*l�B.?~ #��\�����4���C>����F�],���x+9z�>������9sIE��͙���~ӧ��|sb��Q�y��ঽ���d�b�s��*��V��l[��Y��i$-/���-$�ڣ��N�YU�7��_��Y�ڝ�d��*g.�D���g+ `U���8't���+w�#p���@ {����yGP�uIE�c ,�Ԟ{�]�/�o����:��~V�rM�D,�ژx{�?Q�`=�آ@�����Ľ�6�/��|��]2S A��0��ɟ�S��� n�%��X���6�k�����+����!�ɞ�����l���ce �?�����wp]�Z}�����c6�M�\
��z�~Isǣ�DSp_����h�v����X�l)b�|S����kR4�;�v.6���JQp���juɎa U�|��#�s�}�-wD��̫�(���ۋ������>x�,y۷m����C�X�d�m1��C����7#9���u�B
`���m�Y>^S�p��趣���Evtt :v#���F8���
�:F�n+̛��m12oO���D�mk��(���;UHw$��G����%�c�v��[Z��M0#|U_��@���*[�}D�u��#^���D@`p��1����W�0HH�� <�y ^����քm���N�ys�"/7��� X���9�!��U' T��e{K���t�&��c�i�8 ��U(u�]_�(¤I����ӑ��a����Q�@TR�I(1\k����A���$`��w"�O
a�̰�b_~��#��$�1��s�7���������-��	�$r��y�a�Znӑ��T�ޠex�؉l � mx�L�"��xW�9��!�A6&�8��z
挽����rq�/�
ڈ����5��@@@��]��w��ߓ)H=�pUZn�"��|�.�	��罳�u����� �W$��V�y����-S5͠�0

��Z�┭q1�1���g����<&�@�$�&�������E��HT�d��?��e���\���8>����矅Ф���f7~��OG��\X�~A�~0Nz�;�S��^�_}}E��@2/8���~�޾?��bM����7����&�x���;G[g�����Ol<u2��a4o�Le\ڮ$:��?�����D����G�!!CiعY3V$�L���!b���j��<��Wa�����<2�o�'c�O#|�3d���	���A�T�a�,��!��#י������R�=+gM�U_8�lݸ�f|u'�'�,��]�+h�\z5�Q�1Ej;#�{z�S=��U��A����Y����2y��f{\ �E�T�]��%�C�$Zӈ	i5z���������u�Z�vp,�v ?��kMI���    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
q  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�ŗL�e��?�S:/#-l�V�[ڪE�$~��+�̴����K�5[?D��r
Q���2��\�\�
qpw�!w�qpp�}����������g�={�����_���~��x����3�x<N����LK/l'jm��Dݢdh!�9\�q������ct�!��`�/�bG$�|���T�p�C�n�H�87z��}���(t�y�ʆƠ�UZ��,��������/$U�1�2T4�u�uY��AQ&ܤ�-�]��羱�3�3���Y�-Q����b��.W���FŌ{���9�����y} ^�e�[����C?9����-�����Ijd����A7��ډ)W���0�;�Bw�JV�x`�fv��L�[���~�;���j� r_�[����E�� ��]��y=-$2���F-Ne�.�u�W�>���,���~���Uڲ��������=p˗�����S�����'qlo:;���^�������TӅ�b1�S��4���� �}ռ�{��.����|����׈��S��}ܠ��B0 [�h"ջb11M�����I�r�f���(r�h�7_�>��I��������D��	�*N_�?3�+nK�Z�A]|�x=i��اQԚ��<Z�1�?��xw�)R�����=W�(��zJ�A|�����e�T����^|��Q�����B�e 6�@j
16aDy���́�?荀�1 U@?H����i67F��^�0����9�r���3 ��=Aj��0�7:���ro�0E�e�+L0�&��ez,b����Uj1��ZE��@ ���4@244@�����B�6�Z
�B���pqs�
o����Ǹ{XE�y�r����(����N�z�9^��Apx���,����DYzՐ�]
����.:FĢ4�t�8t�'q�P�a�!3!s�-5FyK�>�����9J�{��9�+� j7����s��A��ZTO�E��|�7�B�Z�/b6F[l��!n)�p�j7�� ���*΀�p��^�
q1�,��l�O�'���W>e�+��� 9��T��v �~}���:j����%a�` ��jH� ¿Y����1��ƚs/e z l N)ϴK�|�Ƨڄ�o�;ci��7zzdͳ(��������O��/��wh�Y�f�������'�4���    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
;  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���{PTU��.��*����(G�ɿ��h���5ĀH@��Z(/�ʊ-e�R�͂:>�4LM��U`%b㱬��C���e�',p/2ә��ݳ�����ݳ�,B���� �X,Z��7��R�ɐ|�OYa��L�f��AHr�����p�/q3ψ`�4�����U����T����f��	�����Zr�@P�9�~�C�R �T�s�:nRe^��`��m5�K
�%����ox	j�
�P bP���Dm���մL���M�����X{��otC�Rk^w�{ H~פЬ �����g�%���˫�026��s-8�B0���{��l��Lޗ�>Af�?����7pota�=l�	�k4�I�J��>}����S�İ�&�v�N�0#�<`끓8WG�����<�䕣(s�y@�Ԙ7�����K敡xO�y@<O8��E���"�sX́���F��9��s%������-x�vĮ��Ё4�1�k�廚�
�%p���髳~�*	zEؼ����܀�q�������\��*x�<Cu`Sw�,��F�泍�k�UQU���`����
"HyÏU�W\�uƁ�Z�my-�s���0|��	R����Qu�s�_���W����5@ܗe� -G��-��Vqs�뗍!~�%��@T�>�.%��x0�d$L�p��\���7�`�
<|V��c���yDmm���Q
�-m�����X<Rb;�*ܽ|�澌*
M��u�u@L�R�+C��;0�Å�����?�|%\�=�gA�F��"Ȉ�T1�G��*����)�H���pqu�l�l�u���Po D�."��`P������+<W� '7m{Y��}�P����d�� ؘ^H�3b0(�:��)Z�u��w['g7�ab�O���7�ԑᕾ�y��O5 ���I^f( ���	o,����51�/��N��(U�J����sA�8s��r����`O�u�J �g���vw3F��h�x������x��y�wE�@xr�3(U���q��=!����n�Iq�� �����`?=�Q���P��dv K<����;n�-nY�w#K�����Z���T:8���9���s7>�� ����:~j�*�Nq�?×#��Qx    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
P  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  IDATx�Ŗ{pLWǿK��hR�(�a���LM�Q�iJ�OE<���*��"T}hEDbӄR�JZ�1T��0�?�f�Qb��������{��{z��\�d�n����{�w��;�s��̹G����Ǌ��D���"'�Sw,���0���S䧅��8��%}�EA�t����$ٺh�"��U��2��f�( t���$o���W��`�����`q���	�U��!,�����Mb� �v7����J�5���U
�X��8پl"8/AF�逢���"�����-@U5��'��`я�H����
R��Y�k�q��F����[�+�V)X��()\9	.N���\��i#����?��/�Q���ähջ`<�����ۏa����|��dg����"rv�Q<p�ǯ�����Э�@9�����.�C���9���~Μ�`�7)�dX]^l�{V���Y�}���(��H9�'�]�X�B����'J�S��ݸ�貧��l�WѮ�W������0U��)�63��֥�	�77�
���99�+��a)�N�9��4P�����X�JٌQ	�r_f�!��~F� 	��D�s��w`��_�N;f���εp�>���x���ί�xz)zt�FV�A��0�]��(���V�0k��[;ML`F�⠉�C����i��j�B-vŲ�Qq\�ޯf��\L��;M�`�v7�����|@4}{a@T���=m�m�{���	Z����nr�w��g������؁q%h_@���/�hp��j����,%K7p�ȁ�(@T�9��2~���R�@((�Ё�����X�S`�F6�1��e�K�~1ߘm��A���=����v?��5Ťp�ܠ�@�xh�b��zb�D$0�v�.����Fo����� ���kM7l~���:R@LA L���bֵ�:/���q�����\�n�h�נh����r �������A'�{0T��7?�!�eaa32���:���i�</��_1Cѱٺ��_�X��EX<v�R$d��l�����k��M�$�k���`ݰN���[�����j��ȵ5��C8���87��[f�O9�b�3���<�MJN�s��ۡ�����TK��w-��
C���-�+)/��Պ�3DΝ��`]�p��;9����C弲�*4��C�$n֢���L��C��,m2նƅS�C2l0nT�˲{UYz'�fV;&5E��OT(�]I=����l�Ie��/$��򒳑W}�    IEND�B`�  Left Top� Bitmap
      TApplicationEventsApplicationEventsLeft� Top�    TPF0TPropertiesDialogPropertiesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_propertiesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
PropertiesClientHeight�ClientWidtheColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizee� PixelsPerInch`
TextHeight TButtonOkButtonLeftcTop�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTopWidthZHeightv
ActivePageCommonSheetAnchorsakLeftakTopakRightakBottom TabOrder OnChangePageControlChange 	TTabSheetCommonSheetCaption   Allmänt
DesignSizeRZ  TBevelBevel1LeftTop/Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel1LeftTop:Width,HeightCaptionPlats:ShowAccelChar  
TPathLabelLocationLabelLeftUTop:Width� HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabel	FileLabelLeftUTopWidth� HeightAutoSizeCaption	FileLabelShowAccelChar  TLabelLabel2LeftTopPWidthHeightCaptionStorlek:ShowAccelChar  TLabel	SizeLabelLeftUTopPWidth� HeightAnchorsakLeftakTopakRight AutoSizeCaption	SizeLabelShowAccelChar  TLabelLinksToLabelLabelLeftTopfWidth(HeightCaption   Länkar till:ShowAccelChar  
TPathLabelLinksToLabelLeftUTopfWidth� HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TBevelBevel2LeftTop}Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel3LeftTop� Width;HeightCaption   Filrättigheter:FocusControlRightsFrame  TBevelBevel3LeftTop� Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel4LeftTop� Width!HeightCaptionGrupp:FocusControlGroupComboBox  TLabelLabel5LeftTop� Width$HeightCaption   Ägare:FocusControlOwnerComboBox  TImageFileIconImageLeftTopWidth Height AutoSize	  TBevelRecursiveBevelLeftTop8Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  �TRightsFrameRightsFrameLeftTTop� Width� HeightmTabOrder  	TComboBoxGroupComboBoxLeftUTop� Width� HeightDropDownCount	MaxLength2TabOrderTextGroupComboBoxOnChangeControlChangeOnExitGroupComboBoxExit  	TComboBoxOwnerComboBoxLeftUTop� Width� HeightDropDownCount	MaxLength2TabOrderTextOwnerComboBoxOnChangeControlChangeOnExitOwnerComboBoxExit  	TCheckBoxRecursiveCheckLeftTopBWidth=HeightAnchorsakLeftakTopakRight Caption2   Sätt grupp, ägare och filrättigheter &rekursivtTabOrderOnClickControlChange  TButtonCalculateSizeButtonLeft� TopHWidthPHeightAnchorsakTopakRight Caption	   B&eräknaTabOrder OnClickCalculateSizeButtonClick   	TTabSheetChecksumSheetCaptionKontrollsumma
ImageIndex
DesignSizeRZ  TLabelLabel6LeftTopWidth1HeightCaption
&Algoritm:FocusControlChecksumAlgEdit  	TListViewChecksumViewLeftTop(WidthFHeight)AnchorsakLeftakTopakRightakBottom ColumnsCaptionFilWidthd CaptionKontrollsummaWidthd  ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupChecksumViewContextPopup  	TComboBoxChecksumAlgEditLeftPTop	WidthyHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeChecksumAlgEditChangeOnEnterControlChangeOnExitControlChangeItems.StringsXmd5   TButtonChecksumButtonLeft� TopWidthzHeightAnchorsakTopakRight Caption   B&eräkna kontrollsummaTabOrderOnClickChecksumButtonClick  	TGroupBoxChecksumGroupLeftTop(WidthFHeight)AnchorsakLeftakRightakBottom CaptionKontrollsummaTabOrder
DesignSizeF)  TLabelChecksumUnknownLabelLeft
TopWidthuHeightCaptionChecksumUnknownLabelShowAccelChar  TEditChecksumEditLeft
TopWidth2HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextChecksumEdit     TButton
HelpButtonLeftTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  
TPopupMenuListViewMenuLeftTop� 	TMenuItemCopyCaption&KopieraOnClick	CopyClick    TPF0TRemoteTransferDialogRemoteTransferDialogLeft(Top� HelpType	htKeywordHelpKeywordui_duplicateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRemoteTransferDialogClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight 	TGroupBoxGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize��   TLabelSessionLabelLeft1TopWidthJHeightCaption   Mål&session:FocusControlSessionCombo  TLabelLabel3Left1Top<WidthbHeightCaption   Målfjärr&sökväg:FocusControlDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  	TComboBoxSessionComboLeft1TopWidthXHeightStylecsDropDownListAnchorsakLeftakTopakRight DropDownCount	MaxLength� TabOrder OnChangeSessionComboChange  THistoryComboBoxDirectoryEditLeft1TopLWidthXHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxNotDirectCopyCheckLeft7TopiWidthTHeightAnchorsakLeftakTopakRight Caption#   Dubblera via lokal &temporär kopiaTabOrderOnClickNotDirectCopyCheckClick   TButtonOkButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftPTop� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TRightsFrameRightsFrameLeft Top Width� HeightmTabOrder OnContextPopupFrameContextPopup TLabel
OwnerLabelLeftTopWidth HeightCaption   &ÄgareFocusControlOwnerReadCheck  TLabel
GroupLabelLeftTopWidthHeightCaption&GruppFocusControlGroupReadCheck  TLabelOthersLabelLeftTop,Width!HeightCaptionA&ndraFocusControlOthersReadCheck  TSpeedButtonOthersButtonTagLeft Top)Width8HeightFlat	OnClickRightsButtonsClick  TSpeedButtonGroupButtonTagLeft TopWidth8HeightFlat	OnClickRightsButtonsClick  TSpeedButtonOwnerButtonTagLeft TopWidth8HeightFlat	OnClickRightsButtonsClick  TLabel
OctalLabelLeftTopDWidthHeightCaptionO&ktal:FocusControl	OctalEdit  TGrayedCheckBoxOwnerReadCheckTag Left:TopWidth"HeightHint   LäsCaptionRParentShowHintShowHint	TabOrder OnClickControlChange  TGrayedCheckBoxOwnerWriteCheckTag� Left_TopWidth"HeightHintSkrivCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOwnerExecuteCheckTag@Left� TopWidthHeightHint   Kör/ÖppnaCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupReadCheckTag Left:TopWidth"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupWriteCheckTagLeft_TopWidth!HeightCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupExecuteCheckTagLeft� TopWidthHeightCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersReadCheckTagLeft:Top+Width"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersWriteCheckTagLeft_Top+Width!HeightCaptionWParentShowHintShowHint	TabOrder	OnClickControlChange  TGrayedCheckBoxOthersExecuteCheckTagLeft� Top+WidthHeightCaptionXParentShowHintShowHint	TabOrder
OnClickControlChange  	TCheckBoxDirectoriesXCheckLeftTopYWidth� HeightCaptionAddera &X till katalogerTabOrderOnClickControlChange  TEdit	OctalEditLeft7Top@Width@Height	MaxLengthTabOrderText	OctalEditOnChangeOctalEditChangeOnExitOctalEditExit  TGrayedCheckBoxSetUidCheckTag Left� TopWidthFHeightCaption	   Sätt UIDTabOrderOnClickControlChange  TGrayedCheckBoxSetGIDCheckTag Left� TopWidthFHeightCaption	   Sätt GIDTabOrderOnClickControlChange  TGrayedCheckBoxStickyBitCheckTag Left� Top+WidthFHeightCaption
Sticky bitTabOrderOnClickControlChange  TButtonCloseButtonLeft� TopPWidthKHeightCaption   StängTabOrderVisibleOnClickCloseButtonClick  
TPopupMenuRightsPopupImagesRightsImagesOnPopupRightsPopupPopupLeft� Top; 	TMenuItem	Norights1ActionNoRightsAction  	TMenuItemDefaultrights1ActionDefaultRightsAction  	TMenuItem
Allrights1ActionAllRightsAction  	TMenuItem
Leaveasis1ActionLeaveRightsAsIsAction  	TMenuItemN1Caption-  	TMenuItemCopyAsText1ActionCopyTextAction  	TMenuItemCopyAsOctal1ActionCopyOctalAction  	TMenuItemPaste1ActionPasteAction   TActionListRightsActionsImagesRightsImages	OnExecuteRightsActionsExecuteOnUpdateRightsActionsUpdateLeft� Top TActionNoRightsActionCaption   I&nga rättigheter
ImageIndex ShortCutN@  TActionDefaultRightsActionCaption   Stan&dardrättigheter
ImageIndexShortCutD@  TActionAllRightsActionCaption   &Alla rättigheter
ImageIndexShortCutA@  TActionLeaveRightsAsIsActionCaption   &Lämna oförändradShortCutL@  TActionCopyTextActionCaption&Kopiera som text
ImageIndexShortCutC@  TActionCopyOctalActionCaptionKopiera som &oktalt
ImageIndexShortCutO@  TActionPasteActionCaptionKl&istra in
ImageIndexShortCutV@   TPngImageListRightsImages	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
l  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�}�mH�Q��ϳ��^ܴ�h�--�1]bm�l}�̂�ä~��b�$AIER �EJ��6ɷ�N�d�/ihkj{s�����`��u�r�=���9��s)l�N���%�@��RI�X�YL{n�L&?��/�����O���慃p ��S5E��;�����"z�X�~Fl�d�4�Մdi��X �N��>��<����.�d�������2�k�pb�e��JU!R��tR�#��P1D�g����x�|~�\��W��4[6�ey��8k�`ܩ��t�G���y�P��asa|��=C�*+�H����},�61c�vY���8�Z��@���+���E�ç���l=������y����;B �G��Tub:�9�eg��X��@A{{�����۶=��C��=��g�d��FU����]x�ܫP�����<l?���>O�:���I8���! ��g���+������r�.]�t~��IX �$��1�u+O}��S��� �%<ilB��8�N���!]&A
	�Y^�m�Y������XƧ8��E�+�H	`<_�����1�r!Y*����}��.�!02a�#�L�C�铈_ZD�(
_<^�E���fʤs��{c�~�F�EKp�(�zd��p0����N�Ǒ��$[�#�Z(�P  
����h=�%�s`�S�v;����7�.��$+��,Ҁ    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  mIDATx�cd����x�����@|��?�Jn�/��R���t����{/�iŀ	�q3~u�� S{�F Uď��K���s������L�br@�t���z���{�J�0108�<�u?L������>��;�nU���̷7\�W������e�����t3V��� �� �Mg���1�J(�?��
�ٸ�33�<,���-���{��e�)f�FV�@��3׈7`�s@MP@:p�2��=z����4?�a��`W�>r�x����0;�aƜ�`��g�7����`M9�	s,�`Ӟ��p��-��a��n�1�8w�.B3ԀU[�7�℄-y� :���    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
@  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڅ�HSQǿ�mӵ7*i�$ڔ�b���A��U��0���!B*�!T&%iEP3�DB0J�B݆��sj�j��GK�ԙn2������H���{�9�s�{�RX�Z-���+��L�� :��dh�-����B��9���I��43���Z������c�xh��a�	E��Y8�q7��ڼ5	*� 적CfcM�3Q�9�$�a1�D���/��s����W�N�"#@"��'&�j��
8�ͱ����!�ڪJ��u�������<]�Õ\�^�o���!
|jn��/������>9;���uu����v��?�������? b7Y{W�������*��\kY�ԙl$i��%�����m�HI�ךu�D�1]25�m�/M#~��$I���u(-�D�|ƾ�`��2&W���HwnW��^o�̤'�`4w�U���1.=φ���ͬ���Ao+FRV"ۆ�g�T�,���4���E�8*�O1D��I��`�3������`y��z�s1���������D#-_q� !���i�wvѪH����hX���Ӆ��F[�g��A�a���(E���a�sc�a��t��Ĉ��u))!ʽr�V� Q
!��Q7�����2�A����z"�n�/��&�<��Y��]�����\UɅ    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATxڍ��KSQǿ�%5zQF��A���ڃ= D���>̱��Q�V������Z�(JɈ�ħ��$����L�f�����8E�������p�pB.�>"���+șB5�Y�T��H���)r�����n���"��#y�[T�
8w�	_.E��O݁�l�e�M�Ðo�f���-Iv�a}�Pl4���:�����HG����3�	"���n( ��'t%8Q��I������������"���D�
���B���=}�}���N��`�s8\{$#��;$�������.�������D8|=$�[`碸�:��R�:����g��]������`��&�`��o�5���Ch�h����?�b��ڹJpR��ؐ�nˇ|�$�N��j�:�ZX��q`�:u_9�h���ņ̦$������1�E0�{���[�Dʥ��� 98*����Y� �Хs"��9.����ڇ.����1�Zض��8� �A��i�fv WS�)�_�    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?Cf���X�1&���Ӳþ`��e=��(�g���?�����t���VC��w��?�,����(
>}��p��+���/�c`fu�U���i����,b���/X�t�6�>B�܀��5�gU�0|�1�l�b�7 �u���U�^aX����n/�z�<�K3�}ހHj^�Vu8CL�����S62̪�{	xؙ^���p��+���]�]�6 �i���Ց�Us&�$0T�@x	��y�p��S0�νGs*C��7,�?�&�!�zÄ���)���a��f��_b���æ�g�V�A��[�Vm4�ƃ���>����ˀ�%�n�g����n��y�bj�ex��XAݔ5�^���`��9���EA������YX���m�l]޿�aaC4� FFF����]��%t5�{+���2��s0,j��n@t�/aU���4�c7 �j�"���D��   ,E��d�    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd@���]�����3L߸qm���	����?�#��]@Cmذ6�3��iǪ|��c�~0扌��-���79��Ǘ���cЛ��p���Ƿ�2 `�j�kx0�ۧ�Q$�}K���cL�ݧe�}��2�	�_f��3���.�(G.?dX���1&�_`C�8�1�ytŀ�ߓf�2|��E�ӗ�W�fX���9fVw�N!���_GQ��g2ì�`��Y�b��<��/�e�r�Ê]箂p�gxq�����a���/���;/�_{
f߹���n_AQ��_*��P�������æ�g ���2<�qE�2�4�Y�����j����m�`������E�Y�fWG2T����Hk����l��]>��`[&��(�w_�0���� H��3|z�Er�x9ì�h�����j.
�b��[����a�z��o��vAU�rF\�QU��3 
+�Ed��    IEND�B`�  LefthBitmap
      TPngImageListRightsImages120HeightWidth	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
J  �PNG

   IHDR         ��   	pHYs  �  ��o�d  �IDATxڭ�{L[eƟsiiK/P��ފ��K0��13C�X�e��	n!�q���a̈�4�3A��*"�!8.�1$P`ԁ�����z<��'�%����������y�������bB��x�$�63y�#~V�m����?N�09#�PDS�Q����R��$t]��p���Ź��u-g�
����S,�l��Wg�0-Z켛�$H��� ��}����]NW�ŮV��2�&5���l����58bSr�>��O��.@�Ǧ~�׷l�W`rj�6o�t(62t������B���~\\�X�5,\�Шavv�������s�
P7J��0Ι��w�#�*&"����M-y�zm����=�{FDӘ�7�Zj�ޜ��{0*$���N���wi����"E�1���8���/�m
�{��?QS�$p�A�"AS��hʳ���c@
�L��ھ��F�v�#@N(e�6G�`}U	D"�ϵ{ (�u�ۡ��R����155ni>]��D��t���3LL�,�U�T"F÷��i~=������#o#-e;L�Et��4��g듼�r]Jb|�䴑��6��X{�-xK�h���Q���1 #3OI%P�Z������:�V�3����أM��Cx���X��[����5�߄J!��?�yt�2��+q�������R�9��:��Q�]�"@��Q�x�8W�*��`���b�}�h����۱��%�ml.�������ト�ձ��ə�}�~��k�ʲ��龍����*}g��w�[uc��LE9�XZ�	��q�LZ�W
������E�E����YϳQ	y�|3UxD�����H	�Ŷ�J�UI�l��c���z�C�����^��vW�x)2�¤Cᑸ�I]�l:��KQ�	�R�ߖW8��˾ܽ��GH�����!�p�rte��*Mk�NU��I$[�"�;��C'\\9�{�z��I��9,�^���B����|�'�6��f<��    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
4  �PNG

   IHDR         ��   	pHYs  �  ��o�d  �IDATx�cd�2`�&hl����R�t���Q������~��:sl��4���eab�� #�*,���3��'/����7������2���Ӟ��u���2���o��y�����7��T�D8���_���׏�^��l�A�@{���J:���fx����?�e�9�����1��D>�9)�sW��:}h�:^�m���8�nj��5ܾv��7}`��AR���,�B���2|������mphb��%"(�U������@��+6��j������'����j��6��#BBTx9;+Ã篊��և��^y�b��������Ӈ�.�i�_L�6}"��?noZ2Q��q�W���ceaf��t�faff`ff�,@�(v�$$>��a݂^F���[6�]����a����X��1C,�}�<q%�\8�E����a��`�޾y�pp�.GgWyy���}����ܽA��y������z����-��p��aS3s���"���8��
t����8��^LX��a��`�ݽ}���������AEU��]�ρ�Ν=M����5b�,ư��Y�k�}�ʐ��°f�ZF&V���� ��ѣG	8��JLJ\�a߱�`W�������}a��?���?~l����	��Z.&'%�p��Uh,33��321�����y���4��)ʊ3��x�LX�P�"Р#����Uk72�h;��AlN���������8�  u*$�fՓ    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
/  �PNG

   IHDR         ��   	pHYs  �  ��o�d  �IDATxڭ�kL[e����۸�r)c�V7!��e�vd��1�������:�%3�8���>�]> �]�ܦ��6'�a�B)E(Z�J	�+p���ٙ�!�bⓜ��y���Γ��	��A�/�>3�Q�$��7�,�� X�^�W��x��?�5ڷ4U�� ���w���q�$����B`W�A_�,`zFn�P,�?��$\n�Nxv�u$�&>&J�J����}������i�}��*��9��i����h��l�Q=�)&+ea�8������Q��?�7�	�XT�w>ho1|�ʥ�<OIIJ�������`�o?��\o
L��y).&�V,�9�>�.�W�-U&�ܚb8M=���:}�3���c�5����;�l�W��8U��7)>��9�#c�Z�u���ߞo�(Z�eF �~���w�`���"	;U�"AS���h�ߓ��-]�Y�m�buy�|{��"h���{+K?�@@���U�C�?��;��]���_��=�b#�3^بsM��O=�{�E�ђ����8u�������G<��E�B��f9�}6��=Y�P���[30��D��tc���>�H$������䱣�Z��l������ll�PH��z}�B�mٵ9L"B��,g�������-��D�����[OW'>/+Aq��eb�M�`�I�ζ|:�6/N֬E��}&G���֎E�ҏ
�ua�u�a�ys7J+Kp��;�S�X/}I�����������X���Nͩ�j��E���w-���3?��� �Ἣ
��a0�� ='F�:�d9��.������Yd�o��
�!�������,o��߇xh��1~8�H�Y�k��CN�#h������2N��N;?��e1��3y����Z�M�X�gl���y�U=�[b�w4qˆ`7c~�d�!~؇UO�c����7�����[�{S�1[*Z�-�}������ѯ�����u��)�    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  lIDATxڍ�[OA ���DL0^���41�D� �m)x{h����cK�Eʥ\�TDc����\���KRA��V���m�P����ٝ3_&�e�#��j�0#�⋵�d~D,�3{
�K_��_�Yl�ϧ��[Ol�bA5��Q�V[ 9��Z܌�x����_OB����~�	��4H��B$~��ss�ae=���4tj6`-�c�n� _�-���_���O�|a����X� [16䝬������Y���#���l��� ,Y��}6��Ҁ����c-���$x�c/Y3�+��LOpr�t[�nU�"	z|�g�����ȚYP��~KA�
48��TW���YD��&oĵ�9
����>c�}L��+�$��S�eB�HNL	��Z�i
!��a�d��R�;>~�Ľ�I��`���rB#*� kZ��M��I$S�ChJ2@=�N�	�� ���Z��M-��:��Pg��_4#���U���,Z,��������m�� Mm�[��Y_�r�KB���*�����d\�k���.#���SeY�;q��1�����	��]��A�,{K�z�gLGh#�`f��&�����Ul��Z?ٓ�+}M��r���t�    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  RIDATxڕ��Kq��d���+�'BEzB����\��q���ˡ����Y��?�t�VF�IE�X{4DB(Q\��s�m������>�>p�{qܛ;��[��2���ve�WU̡ؐ��,&������."�%4o>�#��˻T:s^-�7nC5��?��چ���%M~�C��vY��~D���7S��=XL�E4:1��j*e�F�C�j�.����"�]���7͗Y�s��
�
٢���\��]e@}[��V%R�b��{�R�*���Hd���*���5�R��nQ-���1@x��W	�L|×Ν�d<�R���+EPc�#|K4f�8���
����R��2"Xgޮ��ʣ�(���0��������?�d*��E!�j˃�j�`��Y#M��_q ��v������B6��\�:��N`|jZ]8{/>̂Vm�z��L<�;����)
����3'����a�j	TԿ�޲}���o�>�g����0�/	jk������y�ߦ�Ys�Zm�x#p6ȃ*S�Z���Ga�샳��p�y"����`���ʢ��ۏ��Fy���O�+m�������caW�    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  eIDATxڍ��ORa�����n[��^7�~��Ȑ #K7g�j�!���)n��ɚRJYԺ��M�'i6TH S-1L��)����ܼg��>�=;g{	�0 �`s���F�T���C�*amƱ�񣜐�<���:?p8����.�_k�Ծ��=7E�M�������|FTV���l�Qm�R����9�? �g�^�-x��)L=���?Dhb:50�c)�GOK��	}OF��#Ly�P@s���ݑ���^���R1~�QC6R����X\f6c�r�`�����b�*�<t2�=��$��	bK+T�W4�A_mo��	�W��u�`��a75Ԟ^�J�jS��J2��093���U��6�$Y�@t�A�w��Y]���_���D�P �<26���$��<|s;���`��p��	�:����w}h�ʒ`��8|�~*ܱ+j1�{���Y���Xu�I0;W�1g~��",ur�,XA�<5;��EIp����)*�v�f]"Q����k`fo��ڷU��f}14V�/ɲ��݆G%��]�k��kf̺�96T�庒,�X�^���Ҷ��`Ck�YnP^�� Ų�(%� -�j���    IEND�B`�  LeftpBitmap
      TPngImageListRightsImages144HeightWidth	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
N  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d   IDATxڵ�{LSWǿ��qio�Ж�K�7�Ud�B������m�-1B���t_��es�Ő�,f3��ũ��p+U�`T�Z(U�K������(4�Mnι����s��|�9��yVC����XF�K�w��K�3H�VA�{���,Ug/���;�%[��S��h�Tp� �<^X��u�!�auyi�s�gg-Qr���	�b�6kz�^0�s����x=dR	j��
��a���l؀�����ݘfH���v��]{#�ru��ePq(`��Q�I�(5���y�=�-�kX �f�<^�ƿo�{�=�O����1<_3���a����h{�	Ⱥ�19%�r�zz\s�+O�:+�#�F}(��li��l:�9<��༙���Uu0��e�10XPXJ�B�>=�U�̖�j�Ʉ!�f.�G*��)�07t�M�F>+�y��-�odf"^�N-���3���c��w�C؏�A�O�T��H¯R*Yz��aXTV[����-M�GK�����5�@J>?�s��R�>�##Q^yA�T��$�P��T|�����h�f�*��q2:zNL(�w���Y/_����M�� :� @��'�*��d2�����`�|q��O��%���ZDprL6�¾1T*%�-��x��b�7�#8cƌ4M��>-�� v}�,x�GJ+E9������ĩ��_����2�H]��P����y���Z�����H7(=އ0�Y�{83 ����85��׳���]6�@�~��p�r�ݐ�)�:D�#a�;p��+�2��}>\���

3��N�c����\0�h5�S��$��u�V >>�[�����fC���COg���ЪUb[ŵ��^F��{{���غ~���6:e�}L��E�Z$�}�$���GH`��"��m�4m$bH.0cSk���e��O�T�K�mY�X�j���my���4
�,$@ t頪�	��x=N/Ön"�Z��8]�l^�#n���(\4_������ӥB��sc��'����B $�R��t��F#���r��v��?ظr��0N���u���%�c�֣es��e�+�;���������x,I�$��_�q���pu�ӽ��!@A�RZTtU��a1���],x��k�LdҞ�R\����rwx;'�쉋S����e�h�R�������{uT�u��Xo�Kg�"�*&N��WRvE*�F��-T�Yn�������|�e���?ڮ�?fB�(�˵�O5�fe�O    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  |IDATxڵ��OQ���m��
��Z�M0jZ[Q1Fc�|Q��U� ����"�Q� ��$bDE�(�Zli-��B�� D�Q��P����e�eK�K6o�����Λyˁi�T��HB,��&���]@�U?GFϺj�M�Nڸ�$��1�HjV�LX?08��B������i5TWP%�n��ʅs9��a�z��?���@.��>쭯顑_�mz�M� E��h!��J�x>��k/t���>
�C�܏}v1�ZG�#��.�F����=��g��zX�I�Y���tIζΎ����v���x�2%�7Cܸda����>��Гm5h����HP,P��z_�~�5�k*'zii��3�nϓ���lwZ뫗�$���$(B�pvS.������SB�hʝ�^O��~�^C�,KN�׮T�����%�/cH۱�M+`j�t�J�� ty�I����PXV$A ��C�K��zs�mg  gR���,��yPR^��@`�uhM��W/f�� @$�Ҋ�L@��q_����7(�?�RD��B��?(
�jv Ap@�^ �p�Όu>����� �.d"��0J74hqڡ�0��ڳ����Y��um.';@ɹc(E4H�)��5ᔸ��P�w���g@�B����l����P�{�(J��f�p�f >��/�����}g@�R����Fv��S�;e)��k����p";!|��ʁA�0N�#�s� #;@��t\E2��O�Li޻[�6�m��S�8E���=a8�}7Z��H�ol���CE��4N�o�{�dΠ��Cv�3��cY��V���q��%��~lȧ��t�>���9�|?\�ܿ����-/���[U� OєShS���ܤ��k��Px(�m    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
.  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  �IDATxڵ�L�W��_[�wK)�u�Py�'�NG��=�%�l�b��1�9nn�d��,�n3:�,d���屁i�R(����G�R��E��w] "��&_���{���{�s�e�?f�e�+~���,_'b��1���t:/�Gƾ�W^�{j@�W���T�\*��xC$�N�j����F���FMiA���Ĥ�%+�95���ˠ��p#�_��w�ã#��
���Ɵ���}aI8����������]x�����(]$��t�F�l��l�z��:+ 	����T�H���-:�����R�Rʈ�ձ��l���4r�c�$�z1*\���
�źJSqE5���	I�$��9!$\5������gHL{yy��Ru���N��H(j��C�Zߡ)�x"`��27���ru}����LJs�lH���0L�j8��e_?#`C�V��,�x�}`��ap��2s��<2s��#���
��`�[n����:��D���{�2��]� 1�2bk���~Z@`��N'R�������L |��I�L>�9yE� �?���@���B;���X$jW��ȭ)֢�Ô?�����B���Rey���B����h%��@���҅���f=n�TŮ�Y�0F�C/
s��=8�E*Q�B!.T�p��V����ѽ� "b	ۖp���:��}}]�uǙ=|<ίyo5u���"�w�����w�MwW.VQ�5N�x�2���at]X^K����USSգvf��Y,	��U׊ګ�rCv�$@�13}'rl/w1.�h����K���~8t8�mVԷU��.��a��B�A<�)V���#(:S�ن�s�� 	޿��\��k�C������?�bA(��؎�ܭh��Dм�X��Q~��E��� p���-�{?�gl{$M%� cƾm��T�U�n<-/����� ��.�Cx������"�:�1ڃи��P���<0�PX�[�� ~�������ӒGB!&�����@�H��ݥ&Y��C����� S�y{G���Bc�l��d޸�m��s9�o��cW�&�.�,L
����w�L���t�V���?*�Nx@z�43�Uɶaj�7����`��g�!{��POj�1�D]n#��W���/��ٽ���4#g���0�����r�}�06��Uӝg87���t��/�CIj2�,I"3���{sm����:���k��    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
]  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڵ�[H�a��#� �ˠ�(�����n��`
���d�2�67�X-O�ҥ,��ʒ��Q`�T�``�lɜ��;��}}���݅�����������B����b�e��A�Ne�]��� �\1B=��~���>��pz�	Z� �7�C��L�jZ��oo��q��Qfj@Q�Kr;��͎uf-�7Y19�����Hj@����Fcm=4`޴����<�]0��R����8L�caszy6��_+���� �p��	i*����	�\�5&���?�q��[�DS� ����Z���i ���hJ�lh{�T�-��-�a��j��}���}D[zY�V$����S\UWd������ikN�[���`Lc�#}��k=D[��͍�Z#n�e�*�̤(�������i�h���� ��i���F�M#j�d�������Ū��}��t9�H��#Z����;P],���阣�0!�#�CW��V�]e&��n(�:�*L��saN"��yL��y�%	~@J�]������b��a�i�Q�y}Y�_�����{ dZ`Uh�&;��D�=�T݂����7��E*=@�0��t��s�vDDl�I�a(��`TI�i2�ii	bt�p�U���΢����ƞ���S�CH.��U}'zkυ�����;� �>�    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
G  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڵ��OaƟ9�h�I�=p01����`HH5
� J���b]�Tem�B���
�,%����%b�`��*"-��>�Sk�����<���K~CB���<�B�jha����D�	]�����"�2��7���ۯ!A� �ˁ/2�����Y�������DN	4�#��QXp�,�c��&l�����&�G�%�9ј_���146�|�2�?�@��J0 �~����bna�������Bm� �yq�'kz�&/�R�r��G����4�}��h03�>`�>�ƾQ7�c�7��ԝD[$´30�`y�PMk̊�b�:-=�n�Kܺ3E1�ػ{';��;�dy�PM��D�����m�.Iır.��e����,��B5�.'�bi��;���r*�z��^2���J����M�3����t��Z�Lh�e*
�l����y��f�od���㽀�R�ˏ���
��O�B\����e�g2Eh�͸�c����P��$_e �>�^�<�p��e�i��_遾��?@�6m�>�� �.dG� �
��#]��k��N���b���4ߓh:`R��RdƠ���=Qַ�\�.�Tr��VM�_5���i
�4U~*w���V�Uf
$J����GUkF��Dh A�}�62 }���V�    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx���[HSq��ꡐJ�"�+�zм%�nn�t�E�d���L�9M�""�Ι
Y��Ym�S`)����Kj��9�y��t���-<�H/��p�������;gMӠ(
l��	�$u�9'�n���_`a�m�r����6iH��p�d2x*���|�7M�] �)$�Ŭ�-�d��d��B޶.�,Ϋ|VG�G
4�Pk�C�����)�j��1pƋ�&$@??kN\�F^^.�U��9f X�޶v(���l�r
0��s���G�Y6�CcPOh���p2F�e��f5S] �&�2R�0��@����L��C�G$�3��`�_5��K��8��^v`Q�w;�f��bG �>4�ѩ94����N�%��X��(>�~���`�I��Mvݒ���Ң�[�Up)���09������̂$9��-�{#��ƿ�ԥ"��A��������ab���D�[(L	ż~��m6�~���ϐ^�~���w�-闠�Ȁ�
E�[�,��CTހ�k[�U�w���t��0���`"���i<+p�ˁ��� 7�Ͷ4�EB&ou�<6��(�X_ʮv�j��B�͂ѥ	�e�x$����1�i0��*d7�(���yT�!���8;�
���a��k��`��=%�qPϹ6A��Os�Z����B�V�n6��؇]��΢���� nU�2?~��LT�}�#�L|�Z�&�-���	��_�m��i��<�]��r%���wq}�K�m�~����J$    IEND�B`�  LeftxBitmap
      TPngImageListRightsImages192Height Width 	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  _IDATxڽ�{PT�ǿw��} �./5�JŕG�0c�D��a�1f��5mR46@����6��D����F�Ą&����E@v�� �Dy/�d�}ܞ{$�3�{����������.�Y�Z-a���<�����1�Q��F�N��Z�f*�|��>M�Fn#�ē�2N�����쭫,��Q|0M�Z$9B��,��!,X	E�b��{���ن[��ڇ��96�ߕ���G��&�SJ/�|^R��R��Aߠ������B) 	��7�֎o�����W��%�� �S�?����Hnǭ��%&��C�(&�uIh�<DG,�� ����x
�eEO�},פ��STA��K��^�����O�o��r���,q��(\����O"�V�Eq����5��t]Yѿ� Q��u�2`q|t����d|�Gt��J>^�&BA�2P>?!f	[��w�ܮ-=5k����+h��ew��x�����[Zmyq�K\�6<^ɲ����9��|���\ݬ Ԛ�W��>M�O�o�b�^�-;��Fbj�U�b"���۵�Eo�
`�&#�_&y.)�!T׷��p" [g@��I�[R�-ŕF#,6�Q2����f�"��ayL$ʵMp��9�Ң����,��Z7;f��$����Sӳ����x������g�l�9{�x��<�mw_���U���U|>�q��<	r�|&^G�I����Q�5�����lo�=}�@Ȍ�}{�j췀�����G�@����X �5Msx���Y �	x���wvOݥt�����ߪ����*��(�����)�=�]_��3���,.u�����gh��(n�e���{ �_|��oڡb��H�D8YXrg��r>�3��ܺ���,��!Z��-������棽U���b.DFE��LC�:6%�_�����|Y6iǍ�:�:q�3�V�ʏ����X���`hn��g76們��& -���՟YGS�q1Q��%�p���o\� �/� �2	NWN
�9[a�Z8�Tx�>l���I���AoD��A��\�Rt��̬�|�^-_���o`0vt��!yJ�w�䎺�(�KPx��$���&� '����Wq	��4�4("�s��6t��J�@��	$�c=,H���=h0v�}�f�ͦ�`���� $
�����+�,�lh�{9���<��Gϻ���ϐE���Ǡ���Վĥ�P��V� t����ɲWM�,��]/qi��"P����I`S��s��e��4q�zO����G�� �^�6���bE�����v��i�p��6.Xe�y�����*8
�q��9���r�����N���w��y�f�0�;����ېi�ܳlں�o��1 
��@\��pW�����q�*��o�]���=o�y�,�I\�4'��xP���[��?��k/rA��{�*��	�N,�+�L0Y@y�h}%��J$�C@:"'Qlr�&������f7\^ON�՞wO�=;��[`>QRU����3 .'���Z=�
"G��χ*�� *���6B.���Fu� �o�s��ivo�B�`A�������Yє�����/犗�d@���G� H_ˮ&��Q��2D jMf�j]��Z8%���Tcu|a�
u�ϿsLvÍ����!�V������=!	җvr��?��p@s�}�P+�������2X3�Db3#���>��[?�F�2ڕ�`n�lC������B���xR1;I���vf�rz�1z�P%�<Jea��bM���ZF"O!�˿P�Gm�R.Ɨ� ��\�g��6��l`p:�À�����ۖ�֣���2�Ϧ    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  NIDATx�Ŗ{LSw�Ͻ�O��B�樺���Aq��Z�es�,�-�Ȣ�2����m��l�|l��O��ЩZHP�j:��i���`T(���ݯ���Rf�^�ǯMn�s~��9����N1�8T*U)R,�q,��1������0�u���b�^�����-��0�F���0�b ����u�(@ff�@���r}[�(�g(R y�$	�h2|>�������}�\.�7n �2W$OK48��>k&LW$�Ç>�����C��H�$)$��p��?�x��s����N��@�F{���yٙOA�X�[�P��d��ځJD+�E�H��e��L�1 �m]�鯱��W�e���Rk�8U��g�L*���FxЄ������p���H����1(	�r<��J�bo���`��d�4#k�h��	��H`��z��Q�YK_����RI�2g�\h��V��<<����Z��<\�o�ʘ*C���ܯ�-Օ�M���%< BU����	~��\��-� �+�������������a7Wχ�M��t�3�fC���>�v�Y_�	`�r�N��%Y�����C#GQ�o����mb��hiv����	$�7�h�Ǔ��|RcKx����u��X T�����=�����jm��d�%����!�^� ���A?��%X�	��l�.uL ���~s�E�NEo��8pRO�pt"ЭH=q�I&��wKs[Ԛ?�t��e���*�*hr�>�0Ћ3A 5G�i�z#>���+��5��� "��p��z| ���(��T�)?S� 
B�����|�6�I�N�3F�~�^��t��U������{������1 �<)�֙�2m��S_�����2u.-DƮ����!4�����ȞbV��>����H�Q�[
7B�/
���2T	�݆j�}��`�B�� }�UJ?�)I���ņ�=ߺy�ܽK�K$8x����(���������"�'KAW�%��N(-)�웋�`ѳ9 �s��4�1�57qؿ�C���B�z�m��1X�v�_Yy|L��.Y���V��j����"E���)2�H-����pX��k���R�z>F��p�B� �*`2[��--�E�^�SS���U���k^_E��t @�k�-(s���\S�`��XΜ.Sc�#{�t��x���6���b���%n ����ôT��]�&&h���H��	��un �>����S��zGT��(Hb���-���Y7��Y�~r�n���D��>�0p�fUgsE�������o�!A�,�	��;�) 6?Cxw�    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
5  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  �IDATxڽ�T�Uǿ�=`�!�@f�PR��A�%pz����e���-3��QO3�L�:%b�zP�|c�$ۄ��6���ؿ���:m��{������s�{�`�C.��YQD<��Ds�].���uh�j�u�����*8���s��u�xY&9��ȿ�Nv������L��&�Noa�,	
@TDB�%���y[?�&���B�>�`��u6=�����`��4I@X�Q�wc�d"�Ca���`4���� �Cxh0����n0��t��}]�n��K,W�KNM�I�,�����5�#���,�TS;�Id�X�N��F պ8��}������� f��?�g���ӧ�s�Jw
V����64Yw76��<!�60�a�^,�&�M��8Y�'Xv������HN��3<,xr|�$h�`챴�.�M�cG���ǧ�9��ca!A�gL���/tM*����H�9=I `*��8���=��[Z��Hq)e��槂�+I�>>�z��r��ʃ�Q�S2^��ק$_��&.�U�~9|ɩ'I>$̈��Ҋ?�\�V)
?@RJ��1��7�OCye-,Vۧ � �v�D,Z:'�:����l�~A�>3:�Ԍݤ�͚�J���ZQ��@j�+�B�yIq��1Y��<x�����	�9�p�+���|1��`����	���k[sޔ���u��<l�YH��<Ir���t?��A��qLU��ǭol��(�˹�g��>xC:�](��=EnC�0��C����wݕ �1l~��.���_whh��yF=��'K���[ՕlZ�C�����/8���� XBpHy�+@tf����!�lV�.� �,[c��URn+�8������y�݃a�=E
�Ž
�h�ӻ%n�(P�JE����X�`��48 �T����;�V��{�6���K�BR�l�����<�P��vw~�$DR��ڦ;ۺp0��+@�ۯ� I�((*�p�^�Bo�����O�z�8��
�G��%��R*�mϽgv�,VF7V��q4מ���Z�Q$ƾC�G�������m���ٸ�3�r�p����<��"���s��A��̣k�Z�P�K�����`���$$
ƒ����'Fx��Z���|nn.��'y���HY%	C7�$�ů+��������*�S�d0?ؚo��+���/�2���$��{����̇���TA�ݞ��bR��e�h܍��z��G围���+Z�{Ҽ�����˥�Y,;����݆2=@�˔J4�i�GVcZ�L<<�Y��k�\�����iK�B(�aw��+�@_�-����;@�jú7D����x�y����K��OoYa���F�z�݈	����۪�!��nOek���T��Y�v��mD�;�/�I��{�4�
��8�Q�xj���Dta�M�5?hq��V����3�cv��f��hE�NU��+����xI��V-�x`1򛦆�����m��v�OG�;lNT�0@����1VB�W�����{i�v��K�b`m��$$�#�PQU�9l�?�z�]x1�1�g
��h�l��9n�w��FMa����'%p�'���Qp}\%����΁����v,��1&
q���!����4;u���i�;,\j�څ�j�di��Ɔy�j��|g���Dz[��S_F��cb��L��4YXP���~4���tا���y�=qU����d�G��EDy#96���^L����
��͊    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  ]IDATx���P�u��׸
$��J�+�K,����1��<��`�R��%0`c�yFqM��Kq(�
�qbf;��c�	8���ŷ�w����:���w������'��(<�a�><~�I	%�&��E��ٛ>���T�E��w�ȁ���ځ�Ne3��;�E�ȿ@}�i�3�DS�T�:����i;j�@�|�WO��f� �JF�:�&t����7J�	8*ƀ����*I��i�!��րQ��B�����=Rr�������!@{�.���y���8�{Y����Qbn84� ���F\�ُq��J�f�cH>ZC�3٘4��3C�������:ʲ#�����$ّP���!a��Q�	�����δ���I-N�N�l�e/8CIx��.|4�P�W�e�?MI�1��5!��<��⧛]���F�̐H��p5Xv1�J��]�	�r+��
l{= ˖z�ǖN��v|}V�Hv��$'Je��*��9��2!�SHس��M�i�Āro�����p5Xd�F �[F�	��FV�i|�U+�,צ�zTʮ!8h�(��j��z� *CB�1:i/��Y���
����jt���`I�ᶀ�t1U���ra�рe��7*�ի��p5X�Yl��">9�|^P��ր�{�����'��j��x��'y��_�NoĒ%�pcY�mbJ��s�xT��4a-*����	@�YxcP\��,�nnU��T
����)w�Kp����y�ز�=J�F��g�������M��-9Qayx����éñ� ˱'�ή�
���W!4x��tGSs�����
*,�����$���a�����UG�8�eV�J��},��`����!A(!_��O�؎&�-���F �{�P�3G��2J���qB����B�3���;����4�i\�ފd���<Hc��Kb�ߕłu���k��^N^�����8RcwZ��Ic�����&Z4X���[]��O��I/!(���{B��l�{�V��m\�����'>A�m3����M�q0,&� ������]�� w�2��    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx���{L[e�
e1f��8�!�&��،.ˢ�JȨ��-���e�ŹA��T�1���N���had�,�Q'NL�M`�c5iX��Ua=��edI�~=G���~�.����sxE�N�`�a[�����M�V	��z��^ �T�Q���$	N1��š�p�&G�x��J��`>@ֈ��_09�C���I�?�D����>i�j���y2���S4�����ͦԩ$Nր7?>Ii����^?�e��^t�82X��j"k����� �?o�W&`����������x��J[�? X.�8��\?F�ơ/|�=���㔶P��<1 Xz��o.h-��P�� +k�t�"�|�n�>�F��=`[i�`�7�3=�8�7�<�'W�A����(f^��L����
�Q5R:�m=�8�;�w�R�$&����GC����Wfh��
�V�(�r+խX�z6�}�w\�F�ъ�H��wC��g�VX�V�Q��w>2!;�����@~Є}���в��o�
\KS"v� 2����$2��sx$v��&�c��>1 )0Pu�m�UnB݁��.t@YՈ��W��}��\�^���:J�����K�KL@��ǘ��i�4�P�S������5�t[B�|-U["é�K����%��񅭛�i/?׌:�9p,}�0<�Z)��=���\���_���29`={��9�5�
Qx���=s��A��$Hk��S�@�R�p����$��X嫏�*3<�����% 	�^��w�1����_�� �O-h(�
�xD�d������<� Ms;����|.P��,�=@Rh 
,�ۇ��V��&oZ��kn^�"u˥�b��(��e�t��쥻���{�1EU�*d���
I`�4���~<�"N���dOP��8v �= #��(�j�m�nB|\,��HZ���럂�4Wn� 	,>?�~�I�w�O�tg2�㐾�;�$��� 	������*,�N��	B#�L�    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���]LSg�����.�,�l1qqY��%^l7��ksj�����d87��9h�Y�%R�M��-� �u�d�nf#��D\a(��іJ��i{�rL�==t�eOӼ���<�/��H��<�h0�x);{��O�:
y�I�7>���lb���,�*8x�4/�>o;w����:8A���!>)!�!/\!���Ϟ\�Xʝe/���d��lQ����!$,S0�$=D���:������_�ɀy��/%�d�µ�t�Ւ��u� �����;2�8�ƣ��N���:�p����Z�P�4�`�� ����ǻ���l�$�X�A ��v�_�F��a�p.@�)x,�x��p�I�MA��aa�W���m5:�7&�-�
�Q:���0'����P*�5y7�hAW�����Q����v[`Z�Δ�"�! q��]8g}��3|��a��	�
ؔ��}$�}�~��`H�����ˇ���������o;Dof)1=�O��`V쇡\	�������K2^����_@8�{�q�j!�k��������u*�aY������=��q���3� U&��!	hM|FM<lgڻd!¤ϊ�����b����,q��tLJ X2�>?Vc��j��es�x�g|uX-بLÄ�O �R���/��o;eJ3�������̡ 2�po��Z$0@��]�Ō�[��Q�7�lU�8`Cz�o[$���\8�d��Po�
�	�ty@Z*�n����*vo|�T����w��SS0��;�S�� v���p�����r6= �ϣ�h�8`��ݤ	
�b��v�7���f4}VH�����C	`Y1�t�0�����ƥy[������vS �ɸk�P��+��l|��7���=‵۷c�r���9P�ݍI2c���lV��($�nv�G�Ũ�"��8rJ�̳��۩ɑHW����B�.Xb��_ȡWc�i�_�c���FcGy��_"!
�/�O���"��    IEND�B`�  Left� Bitmap
         TPF0�TScpCommanderFormScpCommanderFormLeft� Top HelpType	htKeywordHelpKeywordui_commanderCaptionScpCommanderFormClientHeight�ClientWidth�OldCreateOrder	PixelsPerInch`
TextHeight � 	TSplitterSplitterLeft�Top� WidthHeight*CursorcrSizeWEHintj   |Dra för att ändra proportioner på filpaneler. Dubbelklicka för att bredden på filpanelerna ska lika.ResizeStylersUpdateOnCanResizeSplitterCanResizeOnMovedSplitterMoved  �	TSplitterQueueSplitterTopWidth�  �TTBXDockTopDockWidth�Height� OnContextPopupDockContextPopup TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	OptionstboNoAutoHinttboShowHint 
ShrinkModetbsmWrapStretch	TabOrder TTBXSubmenuItemLocalMenuButtonCaption&LokalHelpKeywordui_commander_menu#localHintC   Ändra layout för lokal panel eller ändra katalog/enhet som visas TTBXItemTBXItem1Action)NonVisualDataModule.LocalChangePathAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXSubmenuItemTBXSubmenuItem2Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemTBXItem2Action&NonVisualDataModule.LocalOpenDirAction  TTBXItemTBXItem3Action/NonVisualDataModule.LocalExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem4Action(NonVisualDataModule.LocalParentDirAction  TTBXItemTBXItem5Action&NonVisualDataModule.LocalRootDirAction  TTBXItemTBXItem6Action&NonVisualDataModule.LocalHomeDirAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem7Action#NonVisualDataModule.LocalBackAction  TTBXItemTBXItem8Action&NonVisualDataModule.LocalForwardAction   TTBXItemTBXItem9Action&NonVisualDataModule.LocalRefreshAction  TTBXItem	TBXItem10Action*NonVisualDataModule.LocalAddBookmarkAction  TTBXItem	TBXItem11Action.NonVisualDataModule.LocalPathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemTBXSubmenuItem3Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i lokal panel TTBXItem	TBXItem12Action,NonVisualDataModule.LocalSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem13Action)NonVisualDataModule.LocalSortByNameAction
GroupIndex	RadioItem	  TTBXItem	TBXItem14Action(NonVisualDataModule.LocalSortByExtAction
GroupIndex	RadioItem	  TTBXItem	TBXItem15Action)NonVisualDataModule.LocalSortByTypeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem16Action,NonVisualDataModule.LocalSortByChangedAction
GroupIndex	RadioItem	  TTBXItem	TBXItem17Action)NonVisualDataModule.LocalSortBySizeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem18Action)NonVisualDataModule.LocalSortByAttrAction
GroupIndex	RadioItem	   TTBXSubmenuItemTBXSubmenuItem4Caption&Visa kolumnerHelpKeywordui_file_panel#selecting_columnsHint$   Välj kolumner som ska visas i panel TTBXItem	TBXItem19Action1NonVisualDataModule.ShowHideLocalNameColumnAction  TTBXItem	TBXItem20Action1NonVisualDataModule.ShowHideLocalSizeColumnAction  TTBXItem	TBXItem21Action1NonVisualDataModule.ShowHideLocalTypeColumnAction  TTBXItem	TBXItem22Action4NonVisualDataModule.ShowHideLocalChangedColumnAction  TTBXItem	TBXItem23Action1NonVisualDataModule.ShowHideLocalAttrColumnAction   TTBXItem
TBXItem221Action%NonVisualDataModule.LocalFilterAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_commander_menu#markHint   Kommandon för markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXSeparatorItemTBXSeparatorItem60  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction  TTBXSeparatorItemTBXSeparatorItem61  TTBXItem
TBXItem212Action'NonVisualDataModule.SelectSameExtAction  TTBXItem
TBXItem213Action)NonVisualDataModule.UnselectSameExtAction   TTBXSubmenuItemTBXSubmenuItem5Caption&FilerHelpKeywordui_commander_menu#filesHint   Kommandon för filoperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem	TBXItem28Action!NonVisualDataModule.NewFileAction  TTBXItem	TBXItem24Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXSubmenuItem	TBXItem26Action%NonVisualDataModule.CurrentEditActionDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem	TBXItem29Action,NonVisualDataModule.CurrentAddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7  TTBXSubmenuItemCurrentCopyItemAction$NonVisualDataModule.RemoteCopyActionDropdownCombo	 TTBXItemCurrentCopyNonQueueItemAction,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItemCurrentCopyQueueItemAction)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem51  TTBXItemCurrentMoveItemAction$NonVisualDataModule.RemoteMoveAction   TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXItem	TBXItem34Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem	TBXItem35Action'NonVisualDataModule.CurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem62  TTBXItem
TBXItem163Action0NonVisualDataModule.CurrentCopyToClipboardAction  TTBXItem	TBXItem36Action NonVisualDataModule.PasteAction2  TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItemCustomCommandsMenuAction,NonVisualDataModule.CustomCommandsFileAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem37Action/NonVisualDataModule.FileListToCommandLineAction  TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action*NonVisualDataModule.FileGenerateUrlAction2   TTBXSubmenuItemTBXSubmenuItem25Caption	   &LåsningHint   Hantera fillås TTBXItem
TBXItem214ActionNonVisualDataModule.LockAction  TTBXItem
TBXItem216Action NonVisualDataModule.UnlockAction   TTBXSeparatorItemTBXSeparatorItem9  TTBXItem	TBXItem41Action+NonVisualDataModule.CurrentPropertiesAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_commander_menu#commandsHintAndra kommandon TTBXItem	TBXItem42Action,NonVisualDataModule.CompareDirectoriesAction  TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItem	TBXItem45Action-NonVisualDataModule.SynchronizeBrowsingAction  TTBXItem
TBXItem210Action)NonVisualDataModule.RemoteFindFilesAction  TTBXSubmenuItemQueueSubmenuItemCaption   K&öHelpKeywordui_queue#manageHint   Kommandon för kölistaOnPopupQueueSubmenuItemPopup TTBXItemQueueEnableItem2Action%NonVisualDataModule.QueueEnableAction  TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#manageHint&   Administrationskommandon för kömassa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction  TTBXItem
TBXItem142Action(NonVisualDataModule.QueueDeleteAllAction  TTBXSeparatorItemTBXSeparatorItem39  TTBXItem
TBXItem134Action,NonVisualDataModule.QueueDeleteAllDoneAction    TTBXSubmenuItemTBXSubmenuItem28Action/NonVisualDataModule.CustomCommandsNonFileAction  TTBXSeparatorItemTBXSeparatorItem13  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem	TBXItem58Action*NonVisualDataModule.CloseApplicationAction   TTBXSubmenuItemTBXSubmenuItem19Caption&SessionHelpKeywordui_commander_menu#sessionHint   Kommandon för session TTBXItem
TBXItem113Action$NonVisualDataModule.NewSessionAction  TTBXItem
TBXItem115Action'NonVisualDataModule.CloseSessionAction2  TTBXItem
TBXItem252Action+NonVisualDataModule.DisconnectSessionAction  TTBXItem
TBXItem253Action*NonVisualDataModule.ReconnectSessionAction  TTBXItem
TBXItem218Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem127Action'NonVisualDataModule.RenameSessionAction  TTBXItem
TBXItem114Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem50  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem
TBXItem135Action-NonVisualDataModule.SessionGenerateUrlAction2  TTBXItem
TBXItem227Action(NonVisualDataModule.ChangePasswordAction  TTBXItem	TBXItem76Action*NonVisualDataModule.PrivateKeyUploadAction  TTBXSeparatorItemTBXSeparatorItem23  TTBXColorItemColorMenuItemAction#NonVisualDataModule.ColorMenuActionColorclNone  TTBXSeparatorItemTBXSeparatorItem29  TTBXSubmenuItemTBXSubmenuItem21Action(NonVisualDataModule.OpenedSessionsAction  TTBXSubmenuItemTBXSubmenuItem231Action$NonVisualDataModule.WorkspacesAction  TTBXItem
TBXItem230Action'NonVisualDataModule.SaveWorkspaceAction  TTBXSeparatorItemTBXSeparatorItem53  TTBXSubmenuItemTBXSubmenuItem20Action(NonVisualDataModule.SavedSessionsAction2   TTBXSubmenuItemTBXSubmenuItem9Caption&AlternativHelpKeywordui_commander_menu#optionsHint)   Ändra layout/inställningar för program TTBXSubmenuItemTBXSubmenuItem10Caption   &VerktygsfältHelpKeywordui_toolbarsHint   Visa/dölj verktygsfält TTBXItem	TBXItem64Action/NonVisualDataModule.CommanderCommandsBandAction  TTBXItem	TBXItem60Action.NonVisualDataModule.CommanderSessionBandAction  TTBXItem	TBXItem62Action2NonVisualDataModule.CommanderPreferencesBandAction  TTBXItem	TBXItem63Action+NonVisualDataModule.CommanderSortBandAction  TTBXItem
TBXItem186Action.NonVisualDataModule.CommanderUpdatesBandAction  TTBXItem
TBXItem188Action/NonVisualDataModule.CommanderTransferBandAction  TTBXItem
TBXItem215Action5NonVisualDataModule.CommanderCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem38  TTBXItem	TBXItem74Action"NonVisualDataModule.ToolBar2Action  TTBXSeparatorItemTBXSeparatorItem47  TTBXItem
TBXItem191Action&NonVisualDataModule.LockToolbarsAction  TTBXItem
TBXItem133Action.NonVisualDataModule.SelectiveToolbarTextAction   TTBXSubmenuItemTBXSubmenuItem11Caption&Lokal panelHelpKeywordui_file_panelHint   Ändra layout för lokal panel TTBXItem	TBXItem65Action3NonVisualDataModule.CommanderLocalHistoryBandAction  TTBXItem	TBXItem66Action6NonVisualDataModule.CommanderLocalNavigationBandAction  TTBXItem	TBXItem59Action0NonVisualDataModule.CommanderLocalFileBandAction  TTBXItem	TBXItem61Action5NonVisualDataModule.CommanderLocalSelectionBandAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem67Action#NonVisualDataModule.LocalTreeAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem68Action(NonVisualDataModule.LocalStatusBarAction   TTBXSubmenuItemTBXSubmenuItem12Caption   F&järrpanelHelpKeywordui_file_panelHint   Ändra layout för fjärrpanel TTBXItem	TBXItem69Action4NonVisualDataModule.CommanderRemoteHistoryBandAction  TTBXItem	TBXItem70Action7NonVisualDataModule.CommanderRemoteNavigationBandAction  TTBXItem
TBXItem136Action1NonVisualDataModule.CommanderRemoteFileBandAction  TTBXItem
TBXItem131Action6NonVisualDataModule.CommanderRemoteSelectionBandAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem	TBXItem72Action)NonVisualDataModule.RemoteStatusBarAction   TTBXSeparatorItemTBXSeparatorItem20  TTBXItemSessionsTabsAction3Action&NonVisualDataModule.SessionsTabsAction  TTBXItem	TBXItem73Action*NonVisualDataModule.CommandLinePanelAction  TTBXItem	TBXItem75Action#NonVisualDataModule.StatusBarAction  TTBXSubmenuItemTBXSubmenuItem14Caption   K&öHelpKeywordui_queueHint   Konfigurera kölista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXItem
TBXItem255Action'NonVisualDataModule.QueueFileListAction  TTBXSeparatorItemTBXSeparatorItem22  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action3NonVisualDataModule.QueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem141Action0NonVisualDataModule.QueueSuspendOnceEmptyAction2  TTBXItem
TBXItem224Action1NonVisualDataModule.QueueShutDownOnceEmptyAction2	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXSeparatorItemTBXSeparatorItem49  TTBXItem	TBXItem82Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemRemoteMenuButtonCaption   F&järrHelpKeywordui_commander_menu#remoteHint=   Ändra layout för fjärrpanel eller ändra katalog som visas TTBXItem	TBXItem83Action*NonVisualDataModule.RemoteChangePathAction  TTBXSeparatorItemTBXSeparatorItem24  TTBXSubmenuItemTBXSubmenuItem15Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem90Action'NonVisualDataModule.RemoteRefreshAction  TTBXItem	TBXItem91Action+NonVisualDataModule.RemoteAddBookmarkAction  TTBXItem	TBXItem92Action/NonVisualDataModule.RemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem27  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i fjärrpanel TTBXItem	TBXItem93Action-NonVisualDataModule.RemoteSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem28  TTBXItem	TBXItem94Action*NonVisualDataModule.RemoteSortByNameAction
GroupIndex	RadioItem	  TTBXItem	TBXItem95Action)NonVisualDataModule.RemoteSortByExtAction
GroupIndex	RadioItem	  TTBXItem
TBXItem193Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem	TBXItem96Action-NonVisualDataModule.RemoteSortByChangedAction
GroupIndex	RadioItem	  TTBXItem	TBXItem97Action*NonVisualDataModule.RemoteSortBySizeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem98Action,NonVisualDataModule.RemoteSortByRightsAction
GroupIndex	RadioItem	  TTBXItem	TBXItem99Action+NonVisualDataModule.RemoteSortByOwnerAction
GroupIndex	RadioItem	  TTBXItem
TBXItem100Action+NonVisualDataModule.RemoteSortByGroupAction
GroupIndex	RadioItem	   TTBXSubmenuItemTBXSubmenuItem17Caption&Visa kolumnerHelpKeywordui_file_panel#selecting_columnsHint$   Välj kolumner som ska visas i panel TTBXItem
TBXItem101Action2NonVisualDataModule.ShowHideRemoteNameColumnAction  TTBXItem
TBXItem102Action2NonVisualDataModule.ShowHideRemoteSizeColumnAction  TTBXItem
TBXItem192Action2NonVisualDataModule.ShowHideRemoteTypeColumnAction  TTBXItem
TBXItem103Action5NonVisualDataModule.ShowHideRemoteChangedColumnAction  TTBXItem
TBXItem104Action4NonVisualDataModule.ShowHideRemoteRightsColumnAction  TTBXItem
TBXItem105Action3NonVisualDataModule.ShowHideRemoteOwnerColumnAction  TTBXItem
TBXItem106Action3NonVisualDataModule.ShowHideRemoteGroupColumnAction  TTBXItem
TBXItem179Action8NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction   TTBXItem
TBXItem220Action&NonVisualDataModule.RemoteFilterAction   TTBXSubmenuItemTBXSubmenuItem22Caption   &HjälpHelpKeywordui_commander_menu#helpHint   Hjälp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXItem
TBXItem217ActionNonVisualDataModule.TipsAction  TTBXSeparatorItemTBXSeparatorItem30  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarPreferencesToolbarLeft Top3Caption   InställningarDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem65  TTBXItem
TBXItem256Action'NonVisualDataModule.QueueFileListAction    TTBXToolbarSessionToolbarLeft TopCaptionSessionDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder  TTBXItem
TBXItem123Action$NonVisualDataModule.NewSessionActionDisplayModenbdmImageAndText  TTBXItem
TBXItem219Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem124Action'NonVisualDataModule.CloseSessionAction2  TTBXItem
TBXItem125Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemTBXSubmenuItem23Action(NonVisualDataModule.SavedSessionsAction2DisplayModenbdmImageAndTextOptionstboDropdownArrow    TTBXToolbarSortToolbarLeft TopMCaptionSorteraDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem148Action+NonVisualDataModule.CurrentSortByTypeAction  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarCommandsToolbarLeft TopgCaption	KommandonDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem154Action,NonVisualDataModule.CompareDirectoriesAction  TTBXItem
TBXItem155Action%NonVisualDataModule.SynchronizeAction  TTBXItem
TBXItem156Action)NonVisualDataModule.FullSynchronizeActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem41  TTBXItem
TBXItem157Action!NonVisualDataModule.ConsoleAction  TTBXItem
TBXItem190ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem42  TTBXItem
TBXItem158Action-NonVisualDataModule.SynchronizeBrowsingAction   TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem1Action)NonVisualDataModule.CheckForUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesActionOptions
tboDefault   TTBXSeparatorItemTBXSeparatorItem46  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft-Top� Caption   ÖverföringsinställningarDockPos,DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXLabelItemTransferSettingsLabelItemCaption   ÖverföringsinställningarMargin  TTBXDropDownItemTransferDropDown	EditWidth� Hint0   Välj förinställda överföringsinställningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelCaption    MarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft+Top� CaptionEgna kommandonDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrderVisible   �TPanelRemotePanelLeft�Top� Width�Height*Constraints.MinHeight� Constraints.MinWidth� ParentColor	TabOrder � 
TPathLabelRemotePathLabelLeft TopOWidth�HeightUnixPath	IndentVerticalAutoSizeVertical	HotTrack	OnGetStatusRemotePathLabelGetStatusOnPathClickRemotePathLabelPathClickOnMaskClickRemotePathLabelMaskClickAutoSizeTransparent
OnDblClickPathLabelDblClick  �	TSplitterRemotePanelSplitterLeft Top� Width�HeightCursorcrSizeNSHinti   Dra för att ändra storlek på katalogträd. Dubbelklicka för att gör höjden på katalogträden lika.AlignalTop  �TTBXStatusBarRemoteStatusBarTopWidth�PanelsFramedSize� StretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint    Klicka för att visa dolda filerMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint,   Klicka för att ändra eller ta bort filtretMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis  OnPanelClickRemoteStatusBarPanelClick  �TPanelRemoteDirPanelLeft Top� Width�Height|Constraints.MinHeightF �TUnixDirViewRemoteDirViewWidth�Height|
NortonLikenlOnOnUpdateStatusBarRemoteDirViewUpdateStatusBar	PathLabelRemotePathLabelAddParentDir	OnDDFileOperationExecuted(RemoteFileControlDDFileOperationExecutedOnHistoryGoDirViewHistoryGoOnPathChangeRemoteDirViewPathChange   �TPanelRemoteDrivePanelTopbWidth�Height-AlignalTopConstraints.MinHeight �TUnixDriveViewRemoteDriveViewWidth�Height-TabStop   TTBXDockRemoteTopDockLeft Top Width�HeightOFixAlign	OnContextPopupDockContextPopup TTBXToolbarRemoteHistoryToolbarLeft TopCaption   FjärrhistorikDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemRemoteBackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemRemoteForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	   TTBXToolbarRemoteNavigationToolbarLeftPTopCaption   FjärrnavigeringDockPosHDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem165Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem
TBXItem166Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem
TBXItem167Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem
TBXItem168Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem37  TTBXItem
TBXItem132Action)NonVisualDataModule.RemoteFindFilesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem44  TTBXItem
TBXItem170Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarRemotePathToolbarLeft Top Caption   Fjärrsökväg
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemRemotePathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXSubmenuItemRemoteOpenDirButtonAction'NonVisualDataModule.RemoteOpenDirActionDropdownCombo	OnPopupRemoteOpenDirButtonPopup  TTBXSubmenuItem
TBXItem229Action&NonVisualDataModule.RemoteFilterActionDropdownCombo	 TTBXItem
TBXItem169Action&NonVisualDataModule.RemoteFilterActionOptions
tboDefault   TTBXSeparatorItemTBXSeparatorItem63  TTBXItem
TBXItem237Action/NonVisualDataModule.FileColorsPreferencesAction    TTBXToolbarRemoteFileToolbarLeftTop5Caption   FjärrfilerDockPosDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItem
TBXItem238Action$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem143Action,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItem
TBXItem200Action)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem59  TTBXItem
TBXItem239Action$NonVisualDataModule.RemoteMoveAction   TTBXSeparatorItemTBXSeparatorItem55  TTBXSubmenuItem
TBXItem242Action$NonVisualDataModule.RemoteEditActionDisplayModenbdmImageAndTextDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem
TBXItem241Action&NonVisualDataModule.RemoteDeleteAction  TTBXItem
TBXItem240Action&NonVisualDataModule.RemoteRenameAction  TTBXItem
TBXItem243Action*NonVisualDataModule.RemotePropertiesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem56  TTBXSubmenuItemRemoteNewSubmenuItemCaption&NyDisplayModenbdmImageAndTextHintSkapa objekt|Skapa nytt objekt
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem247Action'NonVisualDataModule.RemoteNewFileAction  TTBXItem
TBXItem244Action*NonVisualDataModule.RemoteCreateDirAction2  TTBXItem
TBXItem246Action,NonVisualDataModule.RemoteAddEditLinkAction2    TTBXToolbarRemoteSelectionToolbarLeftrTop5Caption   FjärrmarkeringDockPos[DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem138Action&NonVisualDataModule.RemoteSelectAction  TTBXItem
TBXItem139Action(NonVisualDataModule.RemoteUnselectAction  TTBXItem
TBXItem140Action)NonVisualDataModule.RemoteSelectAllAction    TTBXDockRemoteBottomDockLeft TopWidth�Height	FixAlign	PositiondpBottom   �TPanel
QueuePanelTopWidth�HeighttParentColor	TabOrder �
TPathLabel
QueueLabelWidth�  �	TSplitterQueueFileListSplitterTop]Width�  �	TListView
QueueView3Width�Height0TabStop  �TTBXDock	QueueDockWidth�  �	TListViewQueueFileListTop`Width�   �TThemePageControlSessionsPageControlTop� Width�  �TPanel
LocalPanelLeft Top� Width�Height*AlignalLeft
BevelOuterbvNoneConstraints.MinHeight� Constraints.MinWidth� ParentBackgroundParentColor	TabOrder  
TPathLabelLocalPathLabelLeft TopOWidth�HeightIndentVerticalAutoSizeVertical	HotTrack	OnGetStatusLocalPathLabelGetStatusOnPathClickLocalPathLabelPathClickOnMaskClickLocalPathLabelMaskClickAutoSize	PopupMenu#NonVisualDataModule.LocalPanelPopupTransparent
OnDblClickPathLabelDblClick  	TSplitterLocalPanelSplitterLeft Top� Width�HeightCursorcrSizeNSHinti   Dra för att ändra storlek på katalogträd. Dubbelklicka för att gör höjden på katalogträden lika.AlignalTopAutoSnapMinSizeFResizeStylersUpdate  TTBXStatusBarLocalStatusBarLeft TopWidth�HeightPanelsFramedSize� StretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint    Klicka för att visa dolda filerMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint,   Klicka för att ändra eller ta bort filtretMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis  ParentShowHintShowHint	UseSystemFontOnClickLocalStatusBarClickOnPanelClickLocalStatusBarPanelClick  TDirViewLocalDirViewLeft Top� Width�Height|AlignalClientConstraints.MinHeightFDoubleBuffered	FullDrag	HideSelectionParentDoubleBuffered	PopupMenu%NonVisualDataModule.LocalDirViewPopupTabOrder	ViewStylevsReportOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterLocalDirViewEnterOnExitDirViewExit	OnKeyDownDirViewKeyDown
OnKeyPressDirViewKeyPressDirColProperties.ExtVisible	PathLabelLocalPathLabelOnUpdateStatusBarLocalDirViewUpdateStatusBarAddParentDir	OnSelectItemDirViewSelectItemOnLoadedDirViewLoadedOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDTargetHasDropHandler"LocalDirViewDDTargetHasDropHandlerOnDDFileOperationLocalFileControlDDFileOperation
OnExecFileLocalDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayConfirmDeleteUseIconUpdateThread	WatchForChanges	OnFileIconForNameLocalDirViewFileIconForNameOnContextPopupLocalDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnHistoryGoDirViewHistoryGoOnPathChangeLocalDirViewPathChangeOnBusyDirViewBusyOnChangeFocusDirViewChangeFocus  TTBXDockLocalTopDockLeft Top Width�HeightOFixAlign	OnContextPopupDockContextPopup TTBXToolbarLocalHistoryToolbarLeft TopCaptionLokal historikDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemLocalBackButtonAction#NonVisualDataModule.LocalBackActionDropdownCombo	  TTBXSubmenuItemLocalForwardButtonAction&NonVisualDataModule.LocalForwardActionDropdownCombo	   TTBXToolbarLocalNavigationToolbarLeftPTopCaptionLokal navigeringDockPosDDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem159Action(NonVisualDataModule.LocalParentDirAction  TTBXItem
TBXItem160Action&NonVisualDataModule.LocalRootDirAction  TTBXItem
TBXItem161Action&NonVisualDataModule.LocalHomeDirAction  TTBXItem
TBXItem162Action&NonVisualDataModule.LocalRefreshAction  TTBXSeparatorItemTBXSeparatorItem43  TTBXItem
TBXItem164Action#NonVisualDataModule.LocalTreeAction   TTBXToolbarLocalPathToolbarLeft Top Caption   Lokal sökväg
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemLocalPathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex!LocalPathComboBoxAdjustImageIndexOnItemClickLocalPathComboBoxItemClickOnCancelLocalPathComboBoxCancel  TTBXSubmenuItemLocalOpenDirButtonAction&NonVisualDataModule.LocalOpenDirActionDropdownCombo	OnPopupLocalOpenDirButtonPopup  TTBXSubmenuItem
TBXItem228Action%NonVisualDataModule.LocalFilterActionDropdownCombo	 TTBXItem
TBXItem245Action%NonVisualDataModule.LocalFilterAction  TTBXSeparatorItemTBXSeparatorItem64  TTBXItem
TBXItem251Action/NonVisualDataModule.FileColorsPreferencesAction    TTBXToolbarLocalFileToolbarLeft Top5CaptionLokala filerDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItem
TBXItem231Action#NonVisualDataModule.LocalCopyActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem144Action+NonVisualDataModule.LocalCopyNonQueueAction  TTBXItem
TBXItem174Action(NonVisualDataModule.LocalCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem58  TTBXItem
TBXItem232Action#NonVisualDataModule.LocalMoveAction   TTBXSeparatorItemTBXSeparatorItem54  TTBXSubmenuItem
TBXItem235Action#NonVisualDataModule.LocalEditActionDisplayModenbdmImageAndTextDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem
TBXItem234Action%NonVisualDataModule.LocalDeleteAction  TTBXItem
TBXItem233Action%NonVisualDataModule.LocalRenameAction  TTBXItem
TBXItem236Action)NonVisualDataModule.LocalPropertiesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem35  TTBXSubmenuItemLocalNewSubmenuItemCaption&NyDisplayModenbdmImageAndTextHintSkapa objekt|Skapa nytt objekt
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem248Action&NonVisualDataModule.LocalNewFileAction  TTBXItem
TBXItem249Action)NonVisualDataModule.LocalCreateDirAction2  TTBXItem
TBXItem250Action+NonVisualDataModule.LocalAddEditLinkAction2    TTBXToolbarLocalSelectionToolbarLeftaTop5CaptionLokal markeringDockPosIDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem137Action%NonVisualDataModule.LocalSelectAction  TTBXItem	TBXItem32Action'NonVisualDataModule.LocalUnselectAction  TTBXItem	TBXItem30Action(NonVisualDataModule.LocalSelectAllAction    
TDriveViewLocalDriveViewLeft TopbWidth�Height-WatchDirectory	DirViewLocalDirViewOnRefreshDrivesLocalDriveViewRefreshDrivesOnBusyDirViewBusyOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDFileOperationLocalFileControlDDFileOperationAlignalTopConstraints.MinHeightDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedTabOrderTabStopOnEnterLocalDriveViewEnterOnNeedHiddenDirectories#LocalDriveViewNeedHiddenDirectories  TTBXDockLocalBottomDockLeft TopWidth�Height	FixAlign	PositiondpBottom   �TTBXDock
BottomDockLeft Top�Width�Height5FixAlign	PositiondpBottomOnContextPopupDockContextPopup TTBXToolbarToolbar2ToolbarLeft TopCaptionSnabbtangenterDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHintStretch	TabOrder Visible TTBXItem
TBXItem171Action'NonVisualDataModule.CurrentRenameActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem172Action%NonVisualDataModule.CurrentEditActionDisplayModenbdmImageAndTextStretch	  TTBXItemCurrentCopyToolbar2ItemAction$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextStretch	  TTBXItemCurrentMoveToolbar2ItemAction$NonVisualDataModule.RemoteMoveActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem175Action*NonVisualDataModule.CurrentCreateDirActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem176Action'NonVisualDataModule.CurrentDeleteActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem177Action+NonVisualDataModule.CurrentPropertiesActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem178Action*NonVisualDataModule.CloseApplicationActionDisplayModenbdmImageAndText
ImageIndex=Stretch	   TTBXToolbarCommandLineToolbarLeft Top CaptionCommandLineToolbarDockModedmCannotFloatStretch	TabOrderVisibleOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXLabelItemCommandLinePromptLabelCaption
CommandX >Margin  TTBXComboBoxItemCommandLineComboOnBeginEditCommandLineComboBeginEditExtendedAccept	OnPopupCommandLineComboPopup    �TTBXStatusBar	StatusBarLeft Top�Width�ImagesGlyphsModule.SessionImagesPanelsSizedStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndex MaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  ParentShowHint	PopupMenu%NonVisualDataModule.CommanderBarPopupShowHint	UseSystemFontOnPanelDblClickStatusBarPanelDblClick  �	TPanelQueueSeparatorPanelLeft TopWidth�HeightAlignalBottom
BevelEdgesbeBottom 	BevelKindbkFlatTabOrder  �TApplicationEventsApplicationEventsLeftHTop`   TPF0�TScpExplorerFormScpExplorerFormLeft� Top� HelpType	htKeywordHelpKeywordui_explorerActiveControlRemoteDirViewCaptionScpExplorerFormClientHeight�ClientWidthxOldCreateOrder	PixelsPerInch`
TextHeight �	TSplitterQueueSplitterTopLWidthx  �TTBXDockTopDockWidthxHeight� OnContextPopupDockContextPopup TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	OptionstboNoAutoHinttboShowHint 
ShrinkModetbsmWrapStretch	TabOrder  TTBXSubmenuItemTBXSubmenuItem5Caption&FilHelpKeywordui_explorer_menu#fileHintFiloperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135Action!NonVisualDataModule.NewFileAction  TTBXItem
TBXItem136Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem20  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXSubmenuItem	TBXItem26Action$NonVisualDataModule.RemoteEditActionDropdownCombo	OnPopupEditMenuItemPopup  TTBXItemTBXItem4Action,NonVisualDataModule.RemoteAddEditLinkAction2  TTBXSeparatorItemTBXSeparatorItem7  TTBXItem	TBXItem34Action&NonVisualDataModule.RemoteDeleteAction  TTBXItem	TBXItem35Action&NonVisualDataModule.RemoteRenameAction  TTBXItem	TBXItem41Action*NonVisualDataModule.RemotePropertiesAction  TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItem	TBXItem30Action$NonVisualDataModule.RemoteCopyActionDropdownCombo	 TTBXItem
TBXItem156Action,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItem
TBXItem158Action)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem39  TTBXItem	TBXItem32Action$NonVisualDataModule.RemoteMoveAction   TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXSeparatorItemTBXSeparatorItem42  TTBXItem	TBXItem62Action0NonVisualDataModule.CurrentCopyToClipboardAction  TTBXItem	TBXItem36Action NonVisualDataModule.PasteAction2  TTBXSeparatorItemTBXSeparatorItem9  TTBXSubmenuItemCustomCommandsMenuAction,NonVisualDataModule.CustomCommandsFileAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action*NonVisualDataModule.FileGenerateUrlAction2   TTBXSubmenuItemTBXSubmenuItem25Caption	   &LåsningHint   Hantera fillås TTBXItem
TBXItem214ActionNonVisualDataModule.LockAction  TTBXItem
TBXItem216Action NonVisualDataModule.UnlockAction   TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem1Action'NonVisualDataModule.CloseSessionAction2  TTBXItemTBXItem2Action*NonVisualDataModule.CloseApplicationAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_explorer_menu#commandsHintAndra kommandon TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItemTBXItem3Action)NonVisualDataModule.RemoteFindFilesAction  TTBXSubmenuItemQueueSubmenuItemCaption   &KöHelpKeywordui_queue#manageHint   Kommandon för kölistaOnPopupQueueSubmenuItemPopup TTBXItemQueueEnableItem2Action%NonVisualDataModule.QueueEnableAction  TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#manageHint&   Administrationskommandon för kömassa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction  TTBXItem
TBXItem154Action(NonVisualDataModule.QueueDeleteAllAction  TTBXSeparatorItemTBXSeparatorItem35  TTBXItem
TBXItem143Action,NonVisualDataModule.QueueDeleteAllDoneAction    TTBXSubmenuItemTBXSubmenuItem28Action/NonVisualDataModule.CustomCommandsNonFileAction  TTBXSeparatorItemTBXSeparatorItem13  TTBXItemTBXItem5Action+NonVisualDataModule.RemoteAddBookmarkAction  TTBXItemTBXItem6Action/NonVisualDataModule.RemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_explorer_menu#markHint   Kommandon för markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXSeparatorItemTBXSeparatorItem41  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction  TTBXSeparatorItemTBXSeparatorItem61  TTBXItem
TBXItem212Action'NonVisualDataModule.SelectSameExtAction  TTBXItem
TBXItem213Action)NonVisualDataModule.UnselectSameExtAction   TTBXSubmenuItemTBXSubmenuItem19CaptionSessionHelpKeywordui_explorer_menu#sessionHint   Kommandon för session TTBXItem
TBXItem113Action$NonVisualDataModule.NewSessionAction  TTBXItem
TBXItem115Action'NonVisualDataModule.CloseSessionAction2  TTBXItem
TBXItem162Action+NonVisualDataModule.DisconnectSessionAction  TTBXItem
TBXItem163Action*NonVisualDataModule.ReconnectSessionAction  TTBXItem	TBXItem90Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem	TBXItem61Action'NonVisualDataModule.RenameSessionAction  TTBXItem
TBXItem114Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem37  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem
TBXItem144Action-NonVisualDataModule.SessionGenerateUrlAction2  TTBXItem
TBXItem160Action(NonVisualDataModule.ChangePasswordAction  TTBXItem	TBXItem14Action*NonVisualDataModule.PrivateKeyUploadAction  TTBXSeparatorItemTBXSeparatorItem23  TTBXColorItemColorMenuItemAction#NonVisualDataModule.ColorMenuActionColorclNone  TTBXSeparatorItemTBXSeparatorItem29  TTBXSubmenuItemTBXSubmenuItem21Action(NonVisualDataModule.OpenedSessionsAction  TTBXSubmenuItemTBXSubmenuItem231Action$NonVisualDataModule.WorkspacesAction  TTBXItem
TBXItem230Action'NonVisualDataModule.SaveWorkspaceAction  TTBXSeparatorItemTBXSeparatorItem53  TTBXSubmenuItemTBXSubmenuItem20Action(NonVisualDataModule.SavedSessionsAction2   TTBXSubmenuItemTBXSubmenuItem1Caption&VisaHelpKeywordui_explorer_menu#viewHint   Ändra layout för program TTBXSubmenuItemTBXSubmenuItem2Caption   &VerktygsfältHelpKeywordui_toolbarsHint   Visa/dölj verktygsfält TTBXItemTBXItem7Action-NonVisualDataModule.ExplorerAddressBandAction  TTBXItemTBXItem8Action-NonVisualDataModule.ExplorerToolbarBandAction  TTBXItemTBXItem9Action/NonVisualDataModule.ExplorerSelectionBandAction  TTBXItem	TBXItem10Action-NonVisualDataModule.ExplorerSessionBandAction  TTBXItem	TBXItem11Action1NonVisualDataModule.ExplorerPreferencesBandAction  TTBXItem	TBXItem12Action*NonVisualDataModule.ExplorerSortBandAction  TTBXItem	TBXItem82Action-NonVisualDataModule.ExplorerUpdatesBandAction  TTBXItem	TBXItem83Action.NonVisualDataModule.ExplorerTransferBandAction  TTBXItem	TBXItem28Action4NonVisualDataModule.ExplorerCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem	TBXItem92Action&NonVisualDataModule.LockToolbarsAction  TTBXItem
TBXItem140Action.NonVisualDataModule.SelectiveToolbarTextAction   TTBXItemSessionsTabsAction3Action&NonVisualDataModule.SessionsTabsAction  TTBXItem	TBXItem13Action#NonVisualDataModule.StatusBarAction  TTBXSubmenuItemTBXSubmenuItem14Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXItem
TBXItem164Action'NonVisualDataModule.QueueFileListAction  TTBXSeparatorItemTBXSeparatorItem22  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action3NonVisualDataModule.QueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem148Action0NonVisualDataModule.QueueSuspendOnceEmptyAction2  TTBXItem
TBXItem224Action1NonVisualDataModule.QueueShutDownOnceEmptyAction2	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXItem	TBXItem15Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXItem	TBXItem16Action%NonVisualDataModule.CurrentIconAction  TTBXItem	TBXItem17Action*NonVisualDataModule.CurrentSmallIconAction  TTBXItem	TBXItem18Action%NonVisualDataModule.CurrentListAction  TTBXItem	TBXItem19Action'NonVisualDataModule.CurrentReportAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemTBXSubmenuItem15Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem20Action'NonVisualDataModule.RemoteRefreshAction  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i panelen TTBXItem	TBXItem93Action-NonVisualDataModule.RemoteSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem28  TTBXItem	TBXItem94Action*NonVisualDataModule.RemoteSortByNameAction
GroupIndex  TTBXItem	TBXItem95Action)NonVisualDataModule.RemoteSortByExtAction
GroupIndex  TTBXItem
TBXItem132Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem	TBXItem96Action-NonVisualDataModule.RemoteSortByChangedAction
GroupIndex  TTBXItem	TBXItem97Action*NonVisualDataModule.RemoteSortBySizeAction
GroupIndex  TTBXItem	TBXItem98Action,NonVisualDataModule.RemoteSortByRightsAction
GroupIndex  TTBXItem	TBXItem99Action+NonVisualDataModule.RemoteSortByOwnerAction
GroupIndex  TTBXItem
TBXItem100Action+NonVisualDataModule.RemoteSortByGroupAction
GroupIndex   TTBXSubmenuItemTBXSubmenuItem17CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint$   Välj kolumner som ska visas i panel TTBXItem
TBXItem101Action2NonVisualDataModule.ShowHideRemoteNameColumnAction  TTBXItem
TBXItem102Action2NonVisualDataModule.ShowHideRemoteSizeColumnAction  TTBXItem
TBXItem131Action2NonVisualDataModule.ShowHideRemoteTypeColumnAction  TTBXItem
TBXItem103Action5NonVisualDataModule.ShowHideRemoteChangedColumnAction  TTBXItem
TBXItem104Action4NonVisualDataModule.ShowHideRemoteRightsColumnAction  TTBXItem
TBXItem105Action3NonVisualDataModule.ShowHideRemoteOwnerColumnAction  TTBXItem
TBXItem106Action3NonVisualDataModule.ShowHideRemoteGroupColumnAction  TTBXItem	TBXItem76Action8NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction   TTBXItem
TBXItem138Action&NonVisualDataModule.RemoteFilterAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem21Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemTBXSubmenuItem22Caption   &HjälpHelpKeywordui_explorer_menu#helpHint   Hjälp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXItem
TBXItem159ActionNonVisualDataModule.TipsAction  TTBXSeparatorItemTBXSeparatorItem30  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarButtonsToolbarLeft Top4Caption	KommandonDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItem
BackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem23Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem24Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem29Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem	TBXItem37Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem24  TTBXItem
TBXItem139Action)NonVisualDataModule.RemoteFindFilesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem15  TTBXSubmenuItem
TBXItem141Action$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem155Action,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItem
TBXItem157Action)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem38  TTBXItem
TBXItem142Action$NonVisualDataModule.RemoteMoveAction   TTBXSeparatorItemTBXSeparatorItem27  TTBXSubmenuItem	TBXItem42Action$NonVisualDataModule.RemoteEditActionDisplayModenbdmImageAndTextDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem	TBXItem45Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem58Action&NonVisualDataModule.RemoteDeleteAction  TTBXItem	TBXItem59Action*NonVisualDataModule.RemotePropertiesActionDisplayModenbdmImageAndText  TTBXItem	TBXItem60Action&NonVisualDataModule.RemoteRenameAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXSubmenuItemNewSubmenuItemCaption&NyDisplayModenbdmImageAndTextHintSkapa objekt|Skapa nytt objekt
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem247Action'NonVisualDataModule.RemoteNewFileAction  TTBXItem
TBXItem244Action*NonVisualDataModule.RemoteCreateDirAction2  TTBXItem
TBXItem246Action,NonVisualDataModule.RemoteAddEditLinkAction2   TTBXItem	TBXItem63Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem91ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem64Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem65Action)NonVisualDataModule.FullSynchronizeActionDisplayModenbdmImageAndText   TTBXToolbarSelectionToolbarLeft TopNCaption	MarkeringDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem	TBXItem66Action NonVisualDataModule.SelectAction  TTBXItem	TBXItem67Action"NonVisualDataModule.UnselectAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem68Action#NonVisualDataModule.SelectAllAction  TTBXItem	TBXItem69Action)NonVisualDataModule.InvertSelectionAction  TTBXItem	TBXItem70Action(NonVisualDataModule.ClearSelectionAction  TTBXItem
TBXItem134Action*NonVisualDataModule.RestoreSelectionAction   TTBXToolbarSessionToolbarLeft TophCaptionSessionDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem123Action$NonVisualDataModule.NewSessionActionDisplayModenbdmImageAndText  TTBXItem
TBXItem137Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem124Action'NonVisualDataModule.CloseSessionAction2  TTBXItem
TBXItem125Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemTBXSubmenuItem23Action(NonVisualDataModule.SavedSessionsAction2DisplayModenbdmImageAndTextOptionstboDropdownArrow    TTBXToolbarPreferencesToolbarLeft Top� Caption   InställningarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXSubmenuItemTBXSubmenuItem3Action+NonVisualDataModule.CurrentCycleStyleActionDropdownCombo	 TTBXItem	TBXItem72Action%NonVisualDataModule.CurrentIconAction  TTBXItem	TBXItem73Action*NonVisualDataModule.CurrentSmallIconAction  TTBXItem	TBXItem74Action%NonVisualDataModule.CurrentListAction  TTBXItem	TBXItem75Action'NonVisualDataModule.CurrentReportAction   TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem44  TTBXItem
TBXItem165Action'NonVisualDataModule.QueueFileListAction   TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarSortToolbarLeft Top� CaptionSorteraDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem133Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarAddressToolbarLeft TopCaptionAdress
DockableTodpTopdpBottom DockModedmCannotFloatDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHint	PopupMenu&NonVisualDataModule.RemoteAddressPopup	ResizableShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize
OnEndModalAddressToolbarEndModal TTBXLabelItemTBXLabelItem1CaptionAdressMargin  TTBXComboBoxItemUnixPathComboBox	EditWidth� OnAcceptTextUnixPathComboBoxAcceptTextOnBeginEditUnixPathComboBoxBeginEdit	ShowImage	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXItem	TBXItem22Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSubmenuItem
TBXItem229Action&NonVisualDataModule.RemoteFilterActionDropdownCombo	 TTBXItem
TBXItem127Action&NonVisualDataModule.RemoteFilterAction  TTBXSeparatorItemTBXSeparatorItem43  TTBXItem
TBXItem161Action/NonVisualDataModule.FileColorsPreferencesAction    TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem4Action)NonVisualDataModule.CheckForUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesActionOptions
tboDefault   TTBXSeparatorItemTBXSeparatorItem46  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft-Top� Caption   ÖverföringsinställningarDockPos,DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXLabelItemTransferSettingsLabelItemCaption   ÖverföringsinställningarMargin  TTBXDropDownItemTransferDropDown	EditWidth� Hint0   Välj förinställda överföringsinställningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelCaption    MarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft+Top� CaptionEgna kommandonDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder	Visible   �TPanelRemotePanelLeft	Top� WidthfHeightfConstraints.MinHeightdConstraints.MinWidth�  �	TSplitterRemotePanelSplitterHeightGHintW   Dra för att ändra storlek på katalogträd. Dubbelklicka för att dölja katalogträd  �TTBXStatusBarRemoteStatusBarTopPWidthfHeightImagesGlyphsModule.SessionImagesPanelsSize� StretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenterHint    Klicka för att visa dolda filerSizexTag TextTruncationtwEndEllipsis 	AlignmenttaCenterHint,   Klicka för att ändra eller ta bort filtretSizexTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndex MaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  OnPanelClickRemoteStatusBarPanelClickOnPanelDblClickStatusBarPanelDblClick  �TPanelRemoteDirPanelWidth�HeightG �TUnixDirViewRemoteDirViewOnUpdateStatusBarRemoteDirViewUpdateStatusBarOnPathChangeRemoteDirViewPathChange   �TPanelRemoteDrivePanelHeightGConstraints.MinWidth(  TTBXDock
BottomDockLeft TopGWidthfHeight	Color	clBtnFaceFixAlign	PositiondpBottom   �TPanel
QueuePanelTopOWidthx �
TPathLabel
QueueLabelWidthx  �	TSplitterQueueFileListSplitterWidthx  �	TListView
QueueView3Widthx  �TTBXDock	QueueDockWidthx  �	TListViewQueueFileListWidthx   �TThemePageControlSessionsPageControlTop� Widthx  �TTBXDockLeftDockLeft Top� Width	HeightfPositiondpLeft  �TTBXDock	RightDockLeftoTop� Width	HeightfPositiondpRight     TPF0TSelectMaskDialogSelectMaskDialogLeftqTopHelpType	htKeywordHelpKeyword	ui_selectBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSelectXClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	Position
poDesignedOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight 	TGroupBox	MaskGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize��   TLabelLabel3LeftTopWidth/HeightCaption	Fil&mask:FocusControlMaskEdit  TLabelColorFileNamesLabelLeftTopVWidth� Height%AnchorsakLeftakTopakBottom AutoSizeCaption!about.html
index.html
photo.jpgColorclWindowParentColorShowAccelCharTransparentWordWrap	  TLabelColorSizesLabelLeft� TopVWidthKHeight%	AlignmenttaRightJustifyAnchorsakLeftakTopakBottom AutoSizeCaptionColorSizesLabelColorclWindowParentColorShowAccelCharTransparentWordWrap	  TLabelColorPaddingLabelLeft� TopVWidth:Height%	AlignmenttaRightJustifyAnchorsakLeftakTopakRightakBottom AutoSizeColorclWindowParentColorShowAccelCharTransparentWordWrap	  	TCheckBoxApplyToDirectoriesCheckLeftTop?Width� HeightCaption   Tillämpa på &katalogerTabOrder  THistoryComboBoxMaskEditLeftTop$WidthHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder Text*.*OnChangeMaskEditChangeOnExitMaskEditExit  TStaticTextHintTextLeft� Top@WidthiHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	  TButton
MaskButtonLeft1Top"WidthPHeightAnchorsakTopakRight Caption	&RedigeraTabOrderOnClickMaskButtonClick  TButtonColorButtonLeft1TopVWidthPHeightAnchorsakTopakRight Caption   &FärgTabOrderOnClickColorButtonClick   TButtonOKBtnLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftMTop� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeftTTop� WidthKHeightAnchorsakRightakBottom Caption&RensaModalResultTabOrderOnClickClearButtonClick     TPF0TSiteAdvancedDialogSiteAdvancedDialogLeft_Top� HelpType	htKeywordHelpKeywordui_login_advancedBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"   Avancerade webbplatsinställningarClientHeight�ClientWidth1Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnClose	FormCloseOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize1� PixelsPerInch`
TextHeight TPanel	MainPanelLeft Top Width1Height�AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlLeft� Top Width�Height�HelpType	htKeyword
ActivePageEnvironmentSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetEnvironmentSheetTagHelpType	htKeywordHelpKeywordui_login_environmentCaption   Miljö
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxEnvironmentGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption   ServermiljöTabOrder 
DesignSize��   TLabelEOLTypeLabelLeftTopWidth� HeightCaption1   Slut på rad &tecken (om det inte ges av server):FocusControlEOLTypeCombo  TLabelUtfLabelLeftTop,Width� HeightCaption   &UTF-8 kodning på filnamn:FocusControlUtfCombo  TLabelTimeDifferenceLabelLeftTopDWidthTHeightCaptionOffset tidszon:FocusControlTimeDifferenceEdit  TLabelTimeDifferenceHoursLabelLeft� TopDWidthHeightAnchorsakTopakRight CaptiontimmarFocusControlTimeDifferenceEdit  TLabelTimeDifferenceMinutesLabelLeftPTopBWidth%HeightAnchorsakTopakRight CaptionminuterFocusControlTimeDifferenceMinutesEdit  	TComboBoxEOLTypeComboLeft@TopWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrder Items.StringsLFCR/LF   	TComboBoxUtfComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder  TUpDownEditTimeDifferenceEditLeft� Top?WidthEHeight	AlignmenttaRightJustifyMaxValue       �@MinValue       ��Value       ��AnchorsakTopakRight TabOrderOnChange
DataChange  TUpDownEditTimeDifferenceMinutesEditLeftTop?WidthEHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��Value       ��AnchorsakTopakRight TabOrderOnChange
DataChange  	TCheckBoxTimeDifferenceAutoCheckLeft� TopZWidth� HeightCaptionIdentifiera &automatisktTabOrderOnClick
DataChange  	TCheckBoxTrimVMSVersionsCheckLeftTopqWidthqHeightCaptionTrimma VMS-versionsnummerTabOrderOnClick
DataChange   	TGroupBoxDSTModeGroupLeft Top� Width�Height]AnchorsakLeftakTopakRight Caption	SommartidTabOrder
DesignSize�]  TRadioButtonDSTModeUnixCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption7   Justera fjärrtidsstämpel med lokal ko&nvention (Unix)TabOrder OnClick
DataChange  TRadioButtonDSTModeWinCheckLeftTop*WidthqHeightAnchorsakLeftakTopakRight Caption-   Justera fjärrtidsstämpel med &DST (Windows)TabOrderOnClick
DataChange  TRadioButtonDSTModeKeepCheckLeftTopAWidthqHeightAnchorsakLeftakTopakRight Caption    Bevara fjärrtidsstämpel (Unix)TabOrderOnClick
DataChange   	TGroupBox
PuttyGroupLeft Top� Width�HeightbAnchorsakLeftakTopakRight CaptionPuTTYTabOrder
DesignSize�b  TLabelPuttySettingsLabelLeftTopWidthtHeightCaption   &PuTTY terminalinställningar:FocusControlEncryptKeyPasswordEdit  TButtonPuttySettingsButtonLeftTop=Width}HeightAnchorsakTopakRight Caption&Redigera i PuTTY...TabOrderOnClickPuttySettingsButtonClick  TEditPuttySettingsEditLeftTop"WidthrHeight	MaxLength@TabOrder TextPuttySettingsEditOnChange
DataChangeOnExitEncryptKeyEditExit    	TTabSheetDirectoriesSheetTagHelpType	htKeywordHelpKeywordui_login_directoriesCaption	Kataloger
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxDirectoriesGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize��   TLabelLocalDirectoryLabelLeftTopoWidthJHeightCaption&Lokal katalogFocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeftTopBWidthWHeightCaption   F&järrkatalogFocusControlRemoteDirectoryEdit  TLabelLocalDirectoryDescLabelLeftTop� Width� HeightCaptionB   Lokal katalog används inte i det utforskar-liknande gränssnittetShowAccelChar  TDirectoryEditLocalDirectoryEditLeftTop� WidthsHeightAcceptFiles	
DialogText    Välj lokal katalog vid uppstartClickKey@AnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChange
DataChange  TEditRemoteDirectoryEditLeftTopSWidthsHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChange
DataChange  	TCheckBoxUpdateDirectoriesCheckLeftTop*WidthqHeightAnchorsakLeftakTopakRight Caption"   Ko&m ihåg senast använda katalogTabOrder  	TCheckBoxSynchronizeBrowsingCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption   Syn&kronisera bläddringTabOrder    	TGroupBoxDirectoryOptionsGroupLeftTop� Width�HeighttAnchorsakLeftakTopakRight Caption   Alternativ vid kalalogläsningTabOrder
DesignSize�t  	TCheckBoxCacheDirectoriesCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption   Cacha &besökta fjärrkatalogerTabOrder OnClick
DataChange  	TCheckBoxCacheDirectoryChangesCheckLeftTop*Width� HeightAnchorsakLeftakTopakRight Caption   Cacha katalogf&örändringarTabOrderOnClick
DataChange  	TCheckBoxResolveSymlinksCheckLeftTopAWidthqHeightAnchorsakLeftakTopakRight Caption   Slå upp symboliska lä&nkarTabOrder  	TCheckBoxPreserveDirectoryChangesCheckLeft� Top*Width� HeightAnchorsakTopakRight Caption&Permanent cacheTabOrder  	TCheckBoxFollowDirectorySymlinksCheckLeftTopXWidthqHeightAnchorsakLeftakTopakRight Caption(   &Följ symboliska länkar till katalogerTabOrder    	TTabSheetRecycleBinSheetTagHelpType	htKeywordHelpKeywordui_login_recycle_binCaptionPapperskorg
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxRecycleBinGroupLeft TopWidth�HeighttAnchorsakLeftakTopakRight CaptionPapperskorgTabOrder 
DesignSize�t  TLabelRecycleBinPathLabelLeftTopBWidth_HeightCaption   Papp&erskorg på servernFocusControlRecycleBinPathEdit  	TCheckBoxDeleteToRecycleBinCheckLeftTopWidthrHeightAnchorsakLeftakTopakRight Caption6   Flytta borttagna filer på servern till &papperskorgenTabOrder OnClick
DataChange  	TCheckBoxOverwrittenToRecycleBinCheckLeftTop*WidthrHeightAnchorsakLeftakTopakRight CaptionG   Flytta &överskrivna filer på servern till papperskorgen (endast SFTP)TabOrderOnClick
DataChange  TEditRecycleBinPathEditLeftTopSWidthrHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRecycleBinPathEditOnChange
DataChange    	TTabSheetEncryptionSheetTagHelpType	htKeywordHelpKeywordui_login_encryptionCaption
Kryptering
TabVisible
DesignSize�~  	TCheckBoxEncryptFilesCheckLeftTopWidth~HeightAnchorsakLeftakTopakRight Caption&Kryptera filerTabOrder OnClick
DataChange  	TGroupBoxEncryptFilesGroupLeft Top Width�HeightyAnchorsakLeftakTopakRight Caption   KrypteringsinställningarTabOrder TLabelLabel13LeftTopWidthKHeightCaptionKrypterings&nyckelFocusControlEncryptKeyPasswordEdit  TEditEncryptKeyVisibleEditLeftTop"WidthrHeight	MaxLength@TabOrderTextEncryptKeyVisibleEditVisibleOnChange
DataChangeOnExitEncryptKeyEditExit  TPasswordEditEncryptKeyPasswordEditLeftTop"WidthrHeight	MaxLength@TabOrder TextEncryptKeyPasswordEditOnChange
DataChangeOnExitEncryptKeyEditExit  	TCheckBoxShowEncryptionKeyCheckLeftTop=WidthuHeightCaption&Visa nyckelTabOrderOnClickShowEncryptionKeyCheckClick  TButtonGenerateKeyButtonLeftTopTWidthuHeightCaption&Generera nyckelTabOrderOnClickGenerateKeyButtonClick    	TTabSheet	SftpSheetTagHelpType	htKeywordHelpKeywordui_login_sftpCaptionSFTP
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxSFTPBugsGroupBoxLeft ToplWidth�HeightFAnchorsakLeftakTopakRight Caption    Upptäckta buggar i SFTP servrarTabOrder
DesignSize�F  TLabelLabel10LeftTopWidth� HeightCaption;   &Omvänd ordning på symboliska länkar i kommandoargument:FocusControlSFTPBugSymlinkCombo  TLabelLabel36LeftTop,Width� HeightCaption3   Feltolkning av filtidsstä&mplar tidigare än 1970:FocusControlSFTPBugSignedTSCombo  	TComboBoxSFTPBugSymlinkComboLeft@TopWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TComboBoxSFTPBugSignedTSComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TGroupBoxSFTPProtocolGroupLeft TopWidth�Height`AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�`  TLabelLabel34LeftTop,Width� HeightCaption"   Före&drar SFTP protokoll version:FocusControlSFTPMaxVersionCombo  TLabelLabel23LeftTopWidth>HeightCaptionSFTP ser&verFocusControlSftpServerEdit  	TComboBoxSFTPMaxVersionComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderItems.Strings0123456   	TComboBoxSftpServerEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextSftpServerEditOnChange
DataChangeItems.StringsStandard/bin/sftp-serversudo su -c /bin/sftp-server   	TCheckBoxAllowScpFallbackCheckLeftTopDWidthqHeightAnchorsakLeftakTopakRight Caption   Tillåt SCP &fallbackTabOrderOnClick
DataChange    	TTabSheetScpSheetTagHelpType	htKeywordHelpKeywordui_login_scpCaption
SCP/ShellX
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxOtherShellOptionsGroupLeft Top� Width�HeightEAnchorsakLeftakTopakRight Caption   Övriga alternativTabOrder
DesignSize�E  	TCheckBoxLookupUserGroupsCheckLeftTopWidth� HeightAllowGrayed	Caption   Slå upp &användargrupperTabOrder OnClick
DataChange  	TCheckBoxClearAliasesCheckLeftTop*Width� HeightCaptionRensa a&liasTabOrderOnClick
DataChange  	TCheckBoxUnsetNationalVarsCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionRensa &nationella variablerTabOrderOnClick
DataChange  	TCheckBoxScp1CompatibilityCheckLeft� Top*Width� HeightAnchorsakLeftakTopakRight Caption%   Använd scp&2 med scp1 kompatibilitetTabOrderOnClick
DataChange   	TGroupBox
ShellGroupLeft TopWidth�HeightFAnchorsakLeftakTopakRight CaptionSkalTabOrder 
DesignSize�F  TLabelLabel19LeftTopWidthHeightCaptionS&kal:FocusControl	ShellEdit  TLabelLabel20LeftTop,WidthhHeightCaption&Returnera kodvariabel:FocusControlReturnVarEdit  	TComboBox	ShellEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrder Text	ShellEditItems.StringsStandard	/bin/bash/bin/ksh/bin/sh	sudo su -   	TComboBoxReturnVarEditLeft� Top'Width� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextReturnVarEditItems.StringsAutomatisk identifiering?status    	TGroupBoxScpLsOptionsGroupLeft TopTWidth�HeightEAnchorsakLeftakTopakRight CaptionListning av katalogerTabOrder
DesignSize�E  TLabelLabel9LeftTopWidthRHeightCaption   &Kommando för listning:FocusControlListingCommandEdit  	TCheckBoxIgnoreLsWarningsCheckLeftTop*Width� HeightCaptionIgnorera LS &varningarTabOrderOnClick
DataChange  	TCheckBoxSCPLsFullTimeAutoCheckLeft� Top*Width� HeightAnchorsakLeftakTopakRight Caption#   Försök att få &full tidsstämpelTabOrderOnClick
DataChange  	TComboBoxListingCommandEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrder TextListingCommandEditItems.Stringsls -lals -gla     	TTabSheetFtpSheetTagHelpType	htKeywordHelpKeywordui_login_ftpCaptionFTP
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxFtpGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize��   TLabelLabel25LeftTop*WidthgHeightCaption&Kommandon efter inloggning:FocusControlPostLoginCommandsMemo  TLabelFtpListAllLabelLeftTop� Width� HeightCaption%   &Support för listning av dolda filerFocusControlFtpListAllCombo  TLabelLabel24LeftTop|Width� HeightCaption,   Använd &MLSD kommandon för kataloglistningFocusControlFtpUseMlsdCombo  TLabelFtpForcePasvIpLabelLeftTop� Width� HeightCaption+   &Tvinga ip-adress för passiva anslutningarFocusControlFtpForcePasvIpCombo  TLabelFtpAccountLabelLeftTopWidth+HeightCaptionK&onto:FocusControlFtpAccountEdit  TLabelLabel3LeftTop� Width� HeightCaption8   Använd &HOST-kommando för att välja värd på servernFocusControlFtpHostCombo  TMemoPostLoginCommandsMemoLeftTop;WidthqHeight5AnchorsakLeftakTopakRight 
ScrollBars
ssVerticalTabOrder  	TComboBoxFtpListAllComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxFtpForcePasvIpComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxFtpUseMlsdComboLeft@TopwWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  TEditFtpAccountEditLeft� TopWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrder TextFtpAccountEditOnChange
DataChange  	TComboBoxFtpHostComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange    	TTabSheetS3SheetTagHelpType	htKeywordHelpKeywordui_login_s3CaptionS3
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxS3GroupLeft TopWidth�HeightFAnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�F  TLabelLabel27LeftTopWidthHHeightCaption&Standardregion:FocusControlS3DefaultReqionCombo  TLabelS3UrlStyleLabelLeftTop,Width1HeightCaption
&URL-stil:FocusControlS3UrlStyleCombo  	TComboBoxS3DefaultReqionComboLeft� TopWidth� HeightAnchorsakLeftakTopakRight 	MaxLength TabOrder TextS3DefaultRegionComboOnChange
DataChangeItems.Strings
af-south-1	ap-east-1ap-northeast-1ap-northeast-2ap-northeast-3
ap-south-1ap-southeast-1ap-southeast-2ca-central-1
cn-north-1cn-northwest-1eu-central-1
eu-north-1
eu-south-1	eu-west-1	eu-west-2	eu-west-3
me-south-1	sa-east-1	us-east-1	us-east-2us-gov-east-1us-gov-west-1	us-west-1	us-west-2   	TComboBoxS3UrlStyleComboLeft� Top'Width� HeightAutoCompleteStylecsDropDownListAnchorsakLeftakTopakRight 	MaxLength2TabOrderItems.Strings   Virtuell värd   Sökväg    	TGroupBoxS3AuthenticationGroupLeftTopRWidth�Height� AnchorsakLeftakTopakRight CaptionAutentiseringTabOrder
DesignSize��   TLabelLabel5LeftTopWidthIHeightCaption   &Säkerhetstoken:  TMemoS3SessionTokenMemoLeftTop$WidthsHeight]AnchorsakLeftakTopakRightakBottom 	MaxLength'TabOrder OnChange
DataChange	OnKeyDownNoteMemoKeyDown    	TTabSheetWebDavSheetTagHelpType	htKeywordHelpKeywordui_login_webdavCaptionWebDAV
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxWebdavGroupLeft TopWidth�Height.AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�.  	TCheckBoxWebDavLiberalEscapingCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption-&Tolerera icke-kodade specialtecken i filnamnTabOrder OnClick
DataChange    	TTabSheet	ConnSheetTagHelpType	htKeywordHelpKeywordui_login_connectionCaption
Anslutning
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxFtpPingGroupLeft Top� Width�HeightuAnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSize�u  TLabelFtpPingIntervalLabelLeftTopZWidth� HeightCaptionSekunder &mellan keepalivesFocusControlFtpPingIntervalSecEdit  TUpDownEditFtpPingIntervalSecEditLeft� TopUWidthIHeight	AlignmenttaRightJustifyMaxValue       �
@MinValue       ��?	MaxLengthTabOrderOnChange
DataChange  TRadioButtonFtpPingOffButtonLeftTopWidthmHeightAnchorsakLeftakTopakRight Caption&AvTabOrder OnClick
DataChange  TRadioButtonFtpPingNullPacketButtonLeftTop*WidthmHeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketEnabledTabOrderOnClick
DataChange  TRadioButtonFtpPingDummyCommandButtonLeftTopAWidthmHeightAnchorsakLeftakTopakRight Caption#   Kör kommandon för &dummy-protkollTabOrderOnClick
DataChange   	TGroupBoxTimeoutGroupLeft TopPWidth�Height.AnchorsakLeftakTopakRight Caption	TimeouterTabOrder
DesignSize�.  TLabelLabel11LeftTopWidthzHeightCaption   Timeout för se&rversvar:FocusControlTimeoutEdit  TLabelLabel12LeftNTopWidth'HeightAnchorsakTopakRight CaptionsekunderFocusControlTimeoutEdit  TUpDownEditTimeoutEditLeft TopWidthIHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@MinValue       �@AnchorsakTopakRight 	MaxLengthTabOrder OnChange
DataChange   	TGroupBox	PingGroupLeft Top� Width�HeightuAnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSize�u  TLabelPingIntervalLabelLeftTopZWidth� HeightCaptionSekunder &mellan keepalivesFocusControlPingIntervalSecEdit  TUpDownEditPingIntervalSecEditLeft TopUWidthIHeight	AlignmenttaRightJustifyMaxValue       �
@MinValue       ��?AnchorsakTopakRight 	MaxLengthTabOrderOnChange
DataChange  TRadioButtonPingOffButtonLeftTopWidthmHeightAnchorsakLeftakTopakRight CaptionA&vTabOrder OnClick
DataChange  TRadioButtonPingNullPacketButtonLeftTop*WidthmHeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketTabOrderOnClick
DataChange  TRadioButtonPingDummyCommandButtonLeftTopAWidthmHeightAnchorsakLeftakTopakRight Caption%   Kör kommandon för &dummy-protokoll:TabOrderOnClick
DataChange   	TGroupBoxIPvGroupLeft Top� Width�Height.AnchorsakLeftakTopakRight Caption   Version för internetprotokollTabOrder TRadioButtonIPAutoButtonLeftTopWidtheHeightCaptionA&utomatiskTabOrder OnClick
DataChange  TRadioButton
IPv4ButtonLeft|TopWidtheHeightCaptionIPv&4TabOrderOnClick
DataChange  TRadioButton
IPv6ButtonLeft� TopWidtheHeightCaptionIPv&6TabOrderOnClick
DataChange   	TGroupBoxConnectionGroupLeft TopWidth�HeightEAnchorsakLeftakTopakRight Caption
AnslutningTabOrder 
DesignSize�E  	TCheckBoxFtpPasvModeCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption   &Passivt lägeTabOrder OnClick
DataChange  	TCheckBoxBufferSizeCheckLeftTop*WidthqHeightAnchorsakLeftakTopakRight Caption(   Optimera storlek på anslutnings&buffertTabOrderOnClick
DataChange    	TTabSheet
ProxySheetTagHelpType	htKeywordHelpKeywordui_login_proxyCaptionProxy
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxProxyTypeGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight CaptionProxyTabOrder 
DesignSize��   TLabelProxyMethodLabelLeftTopWidth9HeightCaption&Typ av proxy:FocusControlSshProxyMethodCombo  TLabelProxyHostLabelLeftTop)WidthUHeightCaption   Pro&xyns värdnamn:FocusControlProxyHostEdit  TLabelProxyPortLabelLeftTop)Width?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlProxyPortEdit  TLabelProxyUsernameLabelLeftTopUWidth7HeightCaption   &Användarnamn:FocusControlProxyUsernameEdit  TLabelProxyPasswordLabelLeft� TopUWidth2HeightCaption   &Lösenord:FocusControlProxyPasswordEdit  	TComboBoxSshProxyMethodComboLeft� TopWidthnHeightStylecsDropDownListTabOrder OnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTPTelnetLokal   TUpDownEditProxyPortEditLeftTop:WidthbHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChange
DataChange  TEditProxyHostEditLeftTop:Width
HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderTextProxyHostEditOnChange
DataChange  TEditProxyUsernameEditLeftTopfWidth� Height	MaxLengthdTabOrderTextProxyUsernameEditOnChange
DataChange  TPasswordEditProxyPasswordEditLeft� TopfWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextProxyPasswordEditOnChange
DataChange  	TComboBoxFtpProxyMethodComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight DropDownCountTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP
SITE %host!USER %proxyuser, USER %user@%host
OPEN %hostUSER %proxyuser, USER %userUSER %user@%hostUSER %proxyuser@%hostUSER %user@%host %proxyuserUSER %user@%proxyuser@%host   	TComboBoxNeonProxyMethodComboLeft� TopWidthnHeightStylecsDropDownListTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP   TButtonProxyAutodetectButtonLeftTop� WidthdHeightCaption&Automatisk identifieringTabOrderOnClickProxyAutodetectButtonClick   	TGroupBoxProxySettingsGroupLeft Top� Width�Height� AnchorsakLeftakTopakRight Caption   Inställningar proxyTabOrder
DesignSize��   TLabelProxyTelnetCommandLabelLeftTopWidthRHeightCaptionTelnetko&mmando:FocusControlProxyTelnetCommandEdit  TLabelLabel17LeftTopcWidth� HeightCaption-   Låt &DNS-namnuppslagningar göras av proxyn:FocusControlProxyDNSCombo  TLabelProxyLocalCommandLabelLeftTopWidthkHeightCaptionLokalt proxyko&mmando:FocusControlProxyLocalCommandEdit  TEditProxyTelnetCommandEditLeftTop#WidthrHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextProxyTelnetCommandEditOnChange
DataChange  	TCheckBoxProxyLocalhostCheckLeftTopMWidthrHeightAnchorsakLeftakTopakRight Caption(   Låt lokala a&nslutningar gå via proxynTabOrder  	TComboBoxProxyDNSComboLeft� Top^Width� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrderItems.Strings
AutomatiskNejJa   TEditProxyLocalCommandEditLeftTop#WidthHeightAnchorsakLeftakTopakRight TabOrderTextProxyLocalCommandEditOnChange
DataChange  TButtonProxyLocalCommandBrowseButtonLeft,Top!WidthRHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClick"ProxyLocalCommandBrowseButtonClick  TStaticTextProxyTelnetCommandHintTextLeft/Top:WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption   mönsterTabOrderTabStop	  TStaticTextProxyLocalCommandHintTextLeft� Top:WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption   mönsterTabOrderTabStop	    	TTabSheetTunnelSheetTagHelpType	htKeywordHelpKeywordui_login_tunnelCaptionTunnel
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxTunnelSessionGroupLeft Top Width�HeightvAnchorsakLeftakTopakRight Caption    Värd för att sätta upp tunnelTabOrder
DesignSize�v  TLabelLabel6LeftTopWidth7HeightCaption   &Värdnamn:FocusControlTunnelHostNameEdit  TLabelLabel14LeftTopWidth?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlTunnelPortNumberEdit  TLabelLabel15LeftTopDWidth7HeightCaption   &Användarnamn:FocusControlTunnelUserNameEdit  TLabelLabel16Left� TopDWidth2HeightCaption   &Lösenord:FocusControlTunnelPasswordEdit  TEditTunnelHostNameEditLeftTop#Width
HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextTunnelHostNameEditOnChange
DataChange  TEditTunnelUserNameEditLeftTopUWidth� Height	MaxLengthdTabOrderTextTunnelUserNameEditOnChange
DataChange  TPasswordEditTunnelPasswordEditLeft� TopUWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextTunnelPasswordEditOnChange
DataChange  TUpDownEditTunnelPortNumberEditLeftTop#WidthbHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChange
DataChange   	TCheckBoxTunnelCheckLeftTopWidth~HeightAnchorsakLeftakTopakRight CaptionAnslut med SSH-tunnelTabOrder OnClick
DataChange  	TGroupBoxTunnelOptionsGroupLeft Top� Width�Height/AnchorsakLeftakTopakRight Caption   Alternativ för tunnelTabOrder
DesignSize�/  TLabelLabel21LeftTopWidthTHeightCaption&Lokal tunnelport:FocusControlTunnelLocalPortNumberEdit  	TComboBoxTunnelLocalPortNumberEditLeftTopWidthbHeightAutoCompleteAnchorsakTopakRight 	MaxLength2TabOrder TextTunnelLocalPortNumberEditOnChange
DataChangeItems.Strings   Välj automatiskt    	TGroupBoxTunnelAuthenticationParamsGroupLeft Top� Width�HeightDAnchorsakLeftakTopakRight CaptionTunnelautentiseringsparametrarTabOrder
DesignSize�D  TLabelLabel18LeftTopWidthKHeightCaptionPrivat nyc&kelfilFocusControlTunnelPrivateKeyEdit3  TFilenameEditTunnelPrivateKeyEdit3LeftTop#WidthrHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEdit3AfterDialogFilter�PuTTY privata nyckelfiler (*.ppk)|*.ppk|Alla privata nyckelfiler (*.ppk;*.pem;*.key;id_*)|*.ppk;*.pem;*.key;id_*|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrder TextTunnelPrivateKeyEdit3OnChange
DataChange    	TTabSheetSslSheetTagHelpType	htKeywordHelpKeywordui_login_tlsCaptionTLS/SSL
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxSslGroupLeft TopWidth�HeightcAnchorsakLeftakTopakRight CaptionTLS/SSL alternativTabOrder 
DesignSize�c  TLabelLabel1LeftTopWidth{HeightCaption   &Lägsta TLS/SSL-version:FocusControlMinTlsVersionCombo  TLabelLabel2LeftTop,WidthHeightCaption   &Högsta TLS/SSL-version:FocusControlMaxTlsVersionCombo  	TComboBoxMinTlsVersionComboLeft0TopWidthMHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChangeMinTlsVersionComboChangeItems.StringsSSL 3.0TLS 1.0TLS 1.1TLS 1.2TLS 1.3   	TComboBoxMaxTlsVersionComboLeft0Top'WidthMHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChangeMaxTlsVersionComboChangeItems.StringsSSL 3.0TLS 1.0TLS 1.1TLS 1.2TLS 1.3   	TCheckBoxSslSessionReuseCheckLeftTopDWidthmHeightAnchorsakLeftakTopakRight Caption6   Å&teranvänd TLS/SSL-sessionsid för dataanslutningarTabOrderOnClick
DataChange   	TGroupBoxTlsAuthenticationGroupLeft TopqWidth�HeightHAnchorsakLeftakTopakRight CaptionParametrar autentiseringTabOrder
DesignSize�H  TLabelLabel4LeftTopWidthcHeightCaptionKlientcertifikatfil:FocusControlTlsCertificateFileEdit  TFilenameEditTlsCertificateFileEditLeftTop%WidthtHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialog!TlsCertificateFileEditAfterDialogFilteriCertifikat och privata nyckelfiler (*.pfx;*.p12;*.key;*.pem)|*.pfx;*.p12;*.key;*.pem|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj klientcertifikatfilenClickKey@AnchorsakLeftakTopakRight TabOrder TextTlsCertificateFileEditOnChange
DataChange    	TTabSheetAdvancedSheetTagHelpType	htKeywordHelpKeywordui_login_sshCaptionSSH
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxProtocolGroupLeft TopWidth�HeightGAnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�G  TLabelLabel37LeftTop*WidthgHeightCaptionSSH protokollversion:FocusControlSshProtCombo2  	TCheckBoxCompressionCheckLeftTopWidthoHeightAnchorsakLeftakTopakRight Caption   Använd &komprimeringTabOrder OnClick
DataChange  	TComboBoxSshProtCombo2Left/Top%WidthPHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChangeItems.Strings   1 (osäker)2    	TGroupBoxEncryptionGroupLeft TopSWidth�Height� AnchorsakLeftakTopakRight Caption   KrypteringsinställningarTabOrder
DesignSize��   TLabelLabel8LeftTopWidth� HeightCaption$   &Riktlinjer för krypteringschiffer:FocusControlCipherListBox  TListBoxCipherListBoxLeftTop$WidthHeightcAnchorsakLeftakTopakRight DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  	TCheckBoxSsh2LegacyDESCheckLeftTop� WidthoHeightAnchorsakLeftakTopakRight Caption-   Tillåt arvsanvänding av single-&DES i SSH-2TabOrder  TButtonCipherUpButtonLeft/Top$WidthPHeightAnchorsakTopakRight Caption&UppTabOrderOnClickCipherButtonClick  TButtonCipherDownButtonLeft/TopDWidthPHeightAnchorsakTopakRight Caption&NerTabOrderOnClickCipherButtonClick    	TTabSheetKexSheetTagHelpType	htKeywordHelpKeywordui_login_kexCaption
Nyckelbyte
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxKexOptionsGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption%   Alternativ för nyckelbytesalgoritmenTabOrder 
DesignSize��   TLabelLabel28LeftTopWidth|HeightCaption   Ri&ktlinjer för algoritmen:FocusControl
KexListBox  TListBox
KexListBoxLeftTop$WidthHeightYAnchorsakLeftakTopakRight DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  TButtonKexUpButtonLeft/Top$WidthPHeightAnchorsakTopakRight Caption&UppTabOrderOnClickKexButtonClick  TButtonKexDownButtonLeft/TopDWidthPHeightAnchorsakTopakRight Caption&NerTabOrderOnClickKexButtonClick  	TCheckBoxAuthGSSAPIKEXCheckLeftTop� WidthHeightCaption!   Försök med &GSSAPI-nyckelutbyteTabOrderOnClick
DataChange   	TGroupBoxKexReexchangeGroupLeft Top� Width�HeightEAnchorsakLeftakTopakRight Caption(   Alternativ för kontroll av nyckelutbyteTabOrder
DesignSize�E  TLabelLabel31LeftTopWidth� HeightCaption?   Max antal minuter innan nyckeluppdatering (0 ger ingen gräns):Color	clBtnFaceFocusControlRekeyTimeEditParentColor  TLabelLabel32LeftTop,Width� HeightCaption<   Max antal data innan nyckeluppdatering (0 ger ingen gräns):Color	clBtnFaceFocusControlRekeyDataEditParentColor  TUpDownEditRekeyTimeEditLeft/TopWidthPHeight	AlignmenttaRightJustifyMaxValue       �	@AnchorsakTopakRight 	MaxLengthTabOrder OnChange
DataChange  TEditRekeyDataEditLeft/Top'WidthPHeightAnchorsakTopakRight 	MaxLength
TabOrderOnChange
DataChange    	TTabSheet	AuthSheetTagHelpType	htKeywordHelpKeywordui_login_authenticationCaptionAutentisering
ImageIndex

TabVisible
DesignSize�~  	TCheckBoxSshNoUserAuthCheckLeftTopWidth~HeightAnchorsakLeftakTopakRight Caption/   Kringgå autentisering helt och hållet (SSH-2)TabOrder OnClick
DataChange  	TGroupBoxAuthenticationGroupLeft Top Width�HeightuAnchorsakLeftakTopakRight Caption   Alternativ för autentiseringTabOrder
DesignSize�u  	TCheckBoxTryAgentCheckLeftTopWidthuHeightAnchorsakLeftakTopakRight Caption,   Försök använda autentisering med &PageantTabOrder OnClick
DataChange  	TCheckBoxAuthTISCheckLeftTopXWidthuHeightAnchorsakLeftakTopakRight Caption=   Försök använda &TIS eller Kryptokort autentisering (SSH-1)TabOrderOnClick
DataChange  	TCheckBoxAuthKICheckLeftTop*WidthuHeightAnchorsakLeftakTopakRight CaptionA   Försök använda 'tangentbords&interaktiv' autentisering (SSH-2)TabOrderOnClick
DataChange  	TCheckBoxAuthKIPasswordCheckLeft TopAWidthaHeightAnchorsakLeftakTopakRight Caption)   Svara med lösenord vid första &promptenTabOrderOnClick
DataChange   	TGroupBoxAuthenticationParamsGroupLeft Top� Width�HeightxAnchorsakLeftakTopakRight CaptionParametrar autentiseringTabOrder
DesignSize�x  TLabelPrivateKeyLabelLeftTop*WidthKHeightCaptionPrivat nyc&kelfilFocusControlPrivateKeyEdit3  	TCheckBoxAgentFwdCheckLeftTopWidthuHeightAnchorsakLeftakTopakRight Caption   Tillåt agent-vidarebe&fordranTabOrder OnClick
DataChange  TFilenameEditPrivateKeyEdit3LeftTop;WidthtHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEdit3AfterDialogFilter�PuTTY privata nyckelfiler (*.ppk)|*.ppk|Alla privata nyckelfiler (*.ppk;*.pem;*.key;id_*)|*.ppk;*.pem;*.key;id_*|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrderTextPrivateKeyEdit3OnChange
DataChange  TButtonPrivateKeyToolsButtonLeft� TopVWidtheHeightCaption&VerktygTabOrderOnClickPrivateKeyToolsButtonClick  TButtonPrivateKeyViewButtonLeftTopVWidth� HeightCaption&Visa publik nyckelTabOrderOnClickPrivateKeyViewButtonClick   	TGroupBoxGSSAPIGroupLeft TopWidth�HeightGAnchorsakLeftakTopakRight CaptionGSSAPITabOrder
DesignSize�G  	TCheckBoxAuthGSSAPICheck3LeftTopWidthuHeightAnchorsakLeftakTopakRight Caption3   Försök använda GSSAPI/SSPI autentisering (SSH-2)TabOrder OnClickAuthGSSAPICheck3Click  	TCheckBoxGSSAPIFwdTGTCheckLeft Top*WidthaHeightAnchorsakLeftakTopakRight Caption4   Tillåt GSSAPI &vidarbefodra autentiseringsuppgifterTabOrderOnClickAuthGSSAPICheck3Click    	TTabSheet	BugsSheetTagHelpType	htKeywordHelpKeywordui_login_bugsCaptionBuggar
ImageIndex	
TabVisible
DesignSize�~  	TGroupBoxBugsGroupBoxLeft TopWidth�Height!AnchorsakLeftakTopakRight Caption   Upptäcka buggar i SSH-servrarTabOrder 
DesignSize�!  TLabelBugIgnore1LabelLeftTop� Width� HeightCaption(Stannar vid &ignore-meddelanden i SSH-1:FocusControlBugIgnore1Combo  TLabelBugPlainPW1LabelLeftTop� Width� HeightCaption*   &Vägrar all lösenordskamouflage i SSH-1:FocusControlBugPlainPW1Combo  TLabelBugRSA1LabelLeftTopWidth� HeightCaption'Stannar vid &RSA-autentisering i SSH-1:FocusControlBugRSA1Combo  TLabelBugHMAC2LabelLeftTopDWidth� HeightCaption(   Beräkningsfel av H&MAC-nycklar i SSH-2:FocusControlBugHMAC2Combo  TLabelBugDeriveKey2LabelLeftTop\Width� HeightCaption.   Beräkningsf&el av krypteringsnycklar i SSH-2:FocusControlBugDeriveKey2Combo  TLabelBugRSAPad2LabelLeftToptWidth� HeightCaption-   Kräver &utfyllnad av RSA-signaturer i SSH-2:FocusControlBugRSAPad2Combo  TLabelBugPKSessID2LabelLeftTop� Width� HeightCaption1Sessio&ns-id i SSH-2 PK autentisering missbrukas:FocusControlBugPKSessID2Combo  TLabelBugRekey2LabelLeftTop� Width� HeightCaption%   Hanterar SSH-2 nyc&kelutbyte dåligt:FocusControlBugRekey2Combo  TLabelBugMaxPkt2LabelLeftTop� Width� HeightCaption+   Ignorerar SSH-2 ma&ximum för paketstorlek:FocusControlBugMaxPkt2Combo  TLabelBugIgnore2LabelLeftTopWidth� HeightCaption(Stannar vid ignore-meddelanden i SSH-&2:FocusControlBugIgnore2Combo  TLabelBugWinAdjLabelLeftTop,Width� HeightCaption,   Stannar på WinSCP:s SSH-2 'winadj' begäranFocusControlBugWinAdjCombo  	TComboBoxBugIgnore1ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugPlainPW1ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder	OnChange
DataChange  	TComboBoxBugRSA1ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder
OnChange
DataChange  	TComboBoxBugHMAC2ComboLeft@Top?Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugDeriveKey2ComboLeft@TopWWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRSAPad2ComboLeft@TopoWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugPKSessID2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRekey2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugMaxPkt2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugIgnore2ComboLeft@TopWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChange
DataChange  	TComboBoxBugWinAdjComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange    	TTabSheet	NoteSheetHelpType	htKeywordHelpKeywordui_login_noteCaption
Anteckning
ImageIndex
TabVisible
DesignSize�~  	TGroupBox	NoteGroupLeft TopWidth�HeightoAnchorsakLeftakTopakRightakBottom Caption
AnteckningTabOrder 
DesignSize�o  TMemoNoteMemoLeftTopWidthsHeightLAnchorsakLeftakTopakRightakBottom 	MaxLength�TabOrder OnChange
DataChange	OnKeyDownNoteMemoKeyDown     TPanel	LeftPanelLeft Top Width� Height�AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� �  	TTreeViewNavigationTreeLeftTop	Width� Height{AnchorsakLeftakTopakRightakBottom DoubleBuffered	HideSelectionHotTrack	IndentParentDoubleBufferedReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChangeOnCollapsingNavigationTreeCollapsingItems.NodeData
W     6               ����           E n v i r o n m e n t X 6               ����            D i r e c t o r i e s X 6               ����            R e c y c l e   b i n X 4           ��������            E n c r y p t i o n X (               ����            S F T P X &               ����            S C P X &           ��������            F T P X $               ����            S 3 X ,           ��������            W e b D A V X 4               ����           C o n n e c t i o n X *               ����            P r o x y X ,               ����            T u n n e l X &               ����           S S H X 8               ����            K e x   e x c h a n g e X <               ����            A u t h e n t i c a t i o n X (               ����            B u g s X (               ����            N o t e X     TButtonOKBtnLeft3Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonColorButtonLeftTop�WidthRHeightAnchorsakLeftakBottom Caption   &FärgTabOrderOnClickColorButtonClick  
TImageListColorImageListAllocByLeft$Top!Bitmap
&  IL  P   �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5                                                                                                                                                                                                                                         K?5 K?5 K?5 K?5                                                                                                                                                                                                                             dYQ K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                         K?5 s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   @            �                       ��� ��      �      �?      �      �      �      �      �      �      �      �      �      �      �      ��      ��                              
TImageListColorImageList120AllocByHeightWidthLeft� Top!Bitmap
�  IL     �������������BM6       6   (   P                                                                                                                                                                                                                                                                                                                                                                                    bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                         K?5 ��o ��o ��o ��o ��o ��o ��o ��o K?5                                                                                                                                                                                                                                                                                         bXO K?5 K?5 0(" 0(" 0(" 0(" K?5 K?5 bXO                                                                                                                                                                                                                                                                                                     '! '! '! '!                                                                                                                                                                                                                                                                                     qg_ K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 qg_                                                                                                                                                                                                                                                         K?5 ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x )�> )�> ��x K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         oe] K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 oe]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   P            �                       ��� ���         ��         ��         ��         ��         �          �          �          �          �          �          �          �          �          �          �          �          �          ���         ���                                 
TImageListColorImageList144AllocByHeightWidthLeft$TopQBitmap
�%  IL h t   �������������BM6       6   (   `              $                                                                                                                                                                                                                                                                                                                                                                                                                                          bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                 K?5 ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o K?5                                                                                                                                                                                                                                                                                                                                                 K?5 s`R s`R s`R K?5 K?5 K?5 K?5 s`R s`R s`R K?5                                                                                                                                                                                                                                                                                                                                                 bXO K?5 K?5 K?5 B7/ B7/ B7/ B7/ K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                                 0(" 0(" 0(" 0("                                                                                                                                                                                                                                                                                                                                             tjc K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 tjc                                                                                                                                                                                                                                                                                                         K?5 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 )�> )�> NB8 K?5                                                                                                                                                                                                                                                                                                         K?5 QD; ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x QD; K?5                                                                                                                                                                                                                                                                                                         K?5 UG= � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � UG= K?5                                                                                                                                                                                                                                                                                                         K?5 XJ? � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � XJ? K?5                                                                                                                                                                                                                                                                                                         K?5 [MB � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � [MB K?5                                                                                                                                                                                                                                                                                                         K?5 ^PD � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ^PD K?5                                                                                                                                                                                                                                                                                                         K?5 bSG � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � bSG K?5                                                                                                                                                                                                                                                                                                         K?5 eUI � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � eUI K?5                                                                                                                                                                                                                                                                                                         K?5 iXL � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � iXL K?5                                                                                                                                                                                                                                                                                                         K?5 l[N � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � l[N K?5                                                                                                                                                                                                                                                                                                         K?5 o^Q � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � o^Q K?5                                                                                                                                                                                                                                                                                                         K?5 saS � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � saS K?5                                                                                                                                                                                                                                                                                                         K?5 vdV � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � vdV K?5                                                                                                                                                                                                                                                                                                         K?5 yfX �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g yfX K?5                                                                                                                                                                                                                                                                                                         ria OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 ria                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   `                                   ��� ���         � ?         � ?         � ?         � ?         ���         �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          ���         ���                                 
TImageListColorImageList192AllocByHeight Width Left� TopQBitmap
�B  IL ` l     �������������BM6       6   (   �               @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  i_W K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 i_W                                                                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o K?5                                                                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 s`R s`R s`R s`R K?5 K?5 K?5 K?5 K?5 K?5 s`R s`R s`R s`R K?5                                                                                                                                                                                                                                                                                                                                                                                                                                                                 i_W K?5 K?5 K?5 K?5 E:1 E:1 E:1 E:1 E:1 E:1 K?5 K?5 K?5 K?5 i_W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     90( 90( 90( 90( 90( 90(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         -&  -&  -&  -&  -&  -&                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��~ L@6 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 L@6 ���                                                                                                                                                                                                                                                                                                                                                                                                                 L@6 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 L@6                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: )�> )�> )�> PC: K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 RE; ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x RE; K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 TG= � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � TG= K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 WI? � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � WI? K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 YK@ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � YK@ K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 [MB � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � [MB K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 ^OD � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ^OD K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 `QF � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � `QF K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 bSG � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � bSG K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 eUI � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � eUI K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 gWK � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � gWK K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 jYL � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � jYL K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 l[N � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � l[N K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 o]P � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � o]P K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 q_R � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � q_R K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 saS � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � saS K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 ucU � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ucU K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 xeW � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � xeW K?5                                                                                                                                                                                                                                                                                                                                                                                                                 L@6 zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY L@6                                                                                                                                                                                                                                                                                                                                                                                                                 ��} K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 L@6 ��~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         BM>       >   (   �                                    ��� ����            ����            �  �            �  �            �  �            �  �            ���            ���            �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              ����            ����                                    
TPopupMenuPrivateKeyMenuLeft� Top� 	TMenuItemPrivateKeyGenerateItemCaption(&Generera nytt nyckelpar med PuTTYgen...OnClickPrivateKeyGenerateItemClick  	TMenuItemPrivateKeyUploadItemCaption%&Installera publik nyckel i server...OnClickPrivateKeyUploadItemClick    TPF0TSymlinkDialogSymlinkDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_symlinkBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSymlinkDialogClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight 	TGroupBoxSymlinkGroupLeftTopWidth|Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize|�   TLabelFileNameLabelLeftTopWidthSHeightCaption   &Länk/genväg fil:FocusControlFileNameEdit  TLabelLabel1LeftTop@WidthgHeightCaption   &Pekar länk/genväg till:FocusControlPointToEdit  TEditFileNameEditLeftTop WidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  TEditPointToEditLeftTopPWidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxHardLinkCheckLeftTopmWidth� HeightCaption   &Hård länkTabOrderOnClickControlChange   TButtonOkButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft8Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TSynchronizeChecklistDialogSynchronizeChecklistDialogLeft4Top� HelpType	htKeywordHelpKeywordui_synchronize_checklistBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionSynchronization checklist XClientHeight	ClientWidth�Color	clBtnFace
ParentFont		Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               [��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��!Z��                                                                                        ![��?y��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��7s��*e��![��                                                                                        ![��j���8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��*e��![��                                                                                        ![��k���9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��9u��+f��![��                                                                                        ![��k���9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��+f��![��                                                                                        ![��k���:w��:w��:w����������������������������������������������������������������������������������������������������������������������������������:w��:w��:w��+g��![��                                                                                        ![��l���;x��;x��;x����������������������������������������������������������������������������������������������������������������������������������;x��;x��;x��,g��![��                                                                                        ![��l���;y��;y��;y����������������������������������������������������������������������������������������������������������������������������������;y��;y��;y��,g��![��                                                                                        ![��l���<z��<z��<z����������������������������������������������������������������������������������������������������������������������������������<z��<z��<z��,h��![��                                                                                        ![��m���={��={��={��������������������������������������������������SO����\X����������������������������������������������������������������������={��={��={��,h��![��                                                                                        ![��m���=|��=|��=|����������������������������������������������B?��������~w������������������������������������������������������������������=|��=|��=|��,i��![��                                                                                        ![��m���>}��>}��>}������������������������������������������B?����������������������������������������������������������������������������>}��>}��>}��-i��![��                                                                                        ![��m���>~��>~��>~��������������������������������������B?��������������x��������������������������������������������������������������>~��>~��>~��-j��![��                                                                                        ![��m���?��?��?����������������������������������B@������������������������������������������������������������������������������?��?��?��-j��![��                                                                                        ![��n���@���@���@�������������������������������B@����������&&����������y����������������������������������������������������������@���@���@���.j��![��                                                                                        ![��n���@���@���@���������������������������B@����������((������je������������������������������������������������������������������@���@���@���.k��![��                                                                                        ![��n���A���A���A�����������������������B@����������((����������������������y������������������������������������������������������A���A���A���.k��![��                                                                                        ![��o���B���B���B�������������������B@����������((������������������jf��������������������������������������������������������������B���B���B���/l��![��                                                                                        ![��o���B���B���B���������������jf����������((����������������������������������z��������������������������������������������������B���B���B���/l��![��                                                                                        ![��o���C���C���C���������������;9��������((������������������������������jf����������������������������������������������������������C���C���C���/m��![��                                                                                        ![��o���C���C���C�����������������������++�����������������������������������������������{����������������������������������������������C���C���C���/m��![��                                                                                        ![��o���D���D���D�������������������������������������������������������������������jg������������������������������������������������������D���D���D���/m��![��                                                                                        ![��p���E���E���E��������������������������������������������������������������������������������{������������������������������������������E���E���E���0m��![��                                                                                        ![��p���E���E���E�����������������������������������������������������������������������kg��������������������������������������������������E���E���E���0n��![��                                                                                        ![��p���F���F���F������������������������������������������������������������������������������������|��������������������������������������F���F���F���0n��![��                                                                                        ![��q���G���G���G���������������������������������������������������������������������������kh����������������������������������������������G���G���G���1o��![��                                                                                        ![��q���G���G���G����������������������������������������������������������������������������������������}����������������������������������G���G���G���1o��![��                                                                                        ![��q���H���H���H�������������������������������������������������������������������������������ki������������������������������������������H���H���H���1p��![��                                                                                        ![��q���H���H���H��������������������������������������������������������������������������������������������}������������������������������H���H���H���1p��![��                                                                                        ![��r���I���I���I�����������������������������������������������������������������������������������ki��������������������������������������I���I���I���1p��![��                                                                                        ![��r���J���J���J������������������������������������������������������������������������������������������������~��������������������������J���J���J���2q��![��                                                                                        ![��r���J���J���J���������������������������������������������������������������������������������������li����������������������������������J���J���J���2q��![��                                                                                        ![��r���K���K���K��������������������������������������������������������������������������������������������������������������������������K���K���K���2r��![��                                                                                        ![��s���L���L���L�������������������������������������������������������������������������������������������lj������������������������������L���L���L���3r��![��                                                                                        ![��s���L���L���L���������������������������������������������������������������������������������������������������������������������������L���L���L���3r��![��                                                                                        ![��s���M���M���M�����������������������������������������������������������������������������������������������lk��������!"������������������M���M���M���3s��![��                                                                                        ![��s���M���M���M���������������������������������������������������������������������������������������������������������++������������������M���M���M���3s��![��                                                                                        ![��t���N���N���N�������������������������������������������������������������������������������������������������������"#��**����������������������N���N���N���4t��![��                                                                                        ![��t���O���O���O�����������������������������������������������������������������������������������������������������������������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O�����������������������������������������������������������������������������������������������������������������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O�����������������������������������������������������������������������������������������������������������������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O�����������������������������������������������������������������������������������������������������������������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O�����������������������������������������������������������������������������������������������������������������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O���������������������������s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O���������������������������s`R�������������������������������������������������������������������������s`R�������������������������O���O���O���4t��![��                                                                                        ![��t���O���O���O���O���O���O���O���O���O���s`R�������������������������������������������������������������������������s`R�![��O���O���O���O���O���O���O���O���4t��![��                                                                                        ![��t���O���O���O���O���O���O���O���O���O���s`R�������������������������������������������������������������������������s`R�![��O���O���O���O���O���O���O���O���4t��![��                                                                                        ![��t���O���O���O���O���O���O���O���O���O���s`R�������������������������������������������������������������������������s`R�![��O���O���O���O���O���O���O���O���4t��![��                                                                                        ![��t���t���t���t���t���t���t���t���t���t���s`R�������������������������������������������������������������������������s`R�![��t���t���t���t���t���t���t���t���D���![��                                                                                         [��![��![��![��![��![��![��![��![��![��![��s`R�������������������������������������������������������������������������s`R�![��![��![��![��![��![��![��![��![��![�� [��                                                                                                                                    s`R������»���������������������ĺ���ym��ym�Ż�����������������������»�����s`R�                                                                                                                                                                                o^N.s_R�s`Rفob�������������Ƽ��s`R�rXOrXOs`R�ǽ���������������ob�s`R�s_R�o^N.                                                                                                                                                                                            o^N.ubT����������xk�lXN        m[R�zm���������taS�o^N.                                                                                                                                                                                                            s_R����������xk�lXN        m[R�zn���������s_R�                                                                                                                                                                                                                r_R����������þ�s`R�p\Rq^Ls`R��þ���������r_R�                                                                                                                                                                                                                r_Qk�������������Ŀ��xl��zn�����������������r_Pi                                                                                                                                                                                                                ``@s`R���������������������������������s_R�UU+                                                                                                                                                                                                                    lXNs`Qϵ�����������������������r`R�lXN                                                                                                                                                                                                                            UU+r_Qnr_Q�s`R�s`R�r_Q�q^PlUU+                                                                                                                                                                                                                                                                                                                                                                                ����������������������������������    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ����  ?�����  ?�������������������������������������������������������������(   0   `          �%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   [��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![�� [��                                                                ![��@z��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��%_��![��                                                                ![��k���:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��:w��+g��![��                                                                ![��l���;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��,g��![��                                                                ![��l���<y��<y��������������������������������������������������������������������������������������������������<y��<y��,g��![��                                                                ![��l���<{��<{��������������������������������������������������������������������������������������������������<{��<{��,h��![��                                                                ![��m���=|��=|��������������������������������������������������������������������������������������������������=|��=|��,i��![��                                                                ![��m���>}��>}��������������������������������������������������������������������������������������������������>}��>}��-i��![��                                                                ![��m���?~��?~������������������������������������������##��<:��������������������������������������������������?~��?~��-j��![��                                                                ![��m���?��?��������������������������������������������oi����������������������������������������������?��?��-j��![��                                                                ![��n���@���@�����������������������������������������������������������������������������������������@���@���.j��![��                                                                ![��n���A���A�������������������������������������������oj������������������������������������������A���A���.k��![��                                                                ![��o���B���B�����������������������������������kf������������������������������������������������B���B���/l��![��                                                                ![��o���B���B�������������������������������ù������#"������pk��������������������������������������B���B���/l��![��                                                                ![��o���C���C���������������������������ú��������������������������������������������������������C���C���/m��![��                                                                ![��o���D���D���������������!!��������Ļ������������������##������pk����������������������������������D���D���/m��![��                                                                ![��p���E���E���������������98������Ļ����������������������������������������������������������������E���E���0m��![��                                                                ![��p���E���E�������������������������������������������������������##������pl������������������������������E���E���0n��![��                                                                ![��p���F���F���������������������������������������������������������������������������������������������F���F���0o��![��                                                                ![��q���G���G�����������������������������������������������������������##������pm��������������������������G���G���1o��![��                                                                ![��q���H���H���������������������������������������������������������������������������������������������H���H���1p��![��                                                                ![��q���H���H���������������������������������������������������������������##������qn����������������������H���H���1p��![��                                                                ![��r���I���I���������������������������������������������������������������������������������������������I���I���1p��![��                                                                ![��r���J���J�������������������������������������������������������������������##������qo������������������J���J���2q��![��                                                                ![��r���K���K���������������������������������������������������������������������������������������������K���K���2q��![��                                                                ![��r���K���K�����������������������������������������������������������������������##������qo��������������K���K���2r��![��                                                                ![��s���L���L���������������������������������������������������������������������������������������������L���L���3r��![��                                                                ![��s���M���M���������������������������������������������������������������������������#$������tr����������M���M���3s��![��                                                                ![��t���N���N�����������������������������������������������������������������������������������88����������N���N���4s��![��                                                                ![��t���N���N�������������������������������������������������������������������������������RQ����������������N���N���4t��![��                                                                ![��t���O���O���������������������������������������������������������������������������������������������������O���O���4t��![��                                                                ![��t���O���O���������������������������������������������������������������������������������������������������O���O���4t��![��                                                                ![��t���O���O���������������������������������������������������������������������������������������������������O���O���4t��![��                                                                ![��t���O���O�����������������������s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R���������������������O���O���4t��![��                                                                ![��t���O���O�����������������������s`R�������������������������������������������������s`R���������������������O���O���4t��![��                                                                ![��t���O���O���O���O���O���O���O���s`R�������������������������������������������������s`R�<��O���O���O���O���O���O���4t��![��                                                                ![��t���O���O���O���O���O���O���O���s`R�������������������������������������������������s`R�<��O���O���O���O���O���O���4t��![��                                                                ![������t���t���t���t���t���t���t���s`R���|���|���|���|���|���|���|���|���|���|���|���|�s`R�R���t���t���t���t���t���t���D���![��                                                                !Z��![��![��![��![��![��![��![��![��s`R���t��������������m`�taR�taR��m`���������������t�s`R�![��![��![��![��![��![��![��![��!Z��                                                                                                    r^NAr`Q�s`R�{hZ�|i\�s`R�s_R�s_R�s`R�|i\�{hZ�s`R�r`Q�r^NA                                                                                                                                                    q\N$r_Q�r_Q�        s_R�r_Q�q\N$                                                                                                                                                                    s`Q�s_Q�        s_Q�s`Q�                                                                                                                                                                        s_R�s`R�s_Q�s_Q�s`R�s_R�                                                                                                                                                                        UU+s_R�s`R�s`R�s_R�UU+                                                                                                                                                                                                                                                                                    ������  ������  ������  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �    �  �����  �����  ������  �����  �����  ������  (   (   P          @                                                                                                                                                                                                           [��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![�� [��                                                ![��@z��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��+g��%`��![��                                                ![��l���;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��;x��,g��![��                                                ![��l���<y������������������������������������������������������������������������������������������<y��,g��![��                                                ![��l���<{������������������������������������������������������������������������������������������<{��,h��![��                                                ![��m���=|������������������������������������������������������������������������������������������=|��,i��![��                                                ![��m���>}��������������������������������������:8��'&����������������������������������������������>}��-i��![��                                                ![��m���?~����������������������������������('������RN������������������������������������������?~��-j��![��                                                ![��m���?������������������������������('����������ȼ��������������������������������������?��-j��![��                                                ![��n���@���������������������������('������������RN��������������������������������������@���.j��![��                                                ![��n���A�����������������������((������((������������Ƚ����������������������������������A���.k��![��                                                ![��o���B�������������������((������((������������������RO����������������������������������B���/l��![��                                                ![��o���B���������������76������((������������������������ȿ������������������������������B���/l��![��                                                ![��o���C���������������((����((������������������������������RO������������������������������C���/m��![��                                                ![��o���D�������������������������������������������������������������������������������������D���/m��![��                                                ![��p���E�����������������������������������������������������������RP��������������������������E���0m��![��                                                ![��p���E�������������������������������������������������������������������������������������E���0n��![��                                                ![��p���F���������������������������������������������������������������SP����������������������F���0o��![��                                                ![��q���G�������������������������������������������������������������������������������������G���1o��![��                                                ![��q���H�������������������������������������������������������������������SQ������������������H���1p��![��                                                ![��q���H��������������������������������������������������������������� ����������������������H���1p��![��                                                ![��r���I�����������������������������������������������������������������������SQ��������������I���1p��![��                                                ![��r���J������������������������������������������������������������������� ������������������J���2q��![��                                                ![��r���K���������������������������������������������������������������������������SR����������K���2q��![��                                                ![��r���K����������������������������������������������������������������������� ��������������K���2r��![��                                                ![��s���L���������������������������������������������������������������������������==��������������L���3r��![��                                                ![��s���M�������������������������������������������������������������������������������������������M���3s��![��                                                ![��t���N�������������������������������������������������������������������������������������������N���4s��![��                                                ![��t���N�������������������������������������������������������������������������������������������N���4t��![��                                                ![��t���O�����������������������s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R���������������������O���4t��![��                                                ![��t���O���O���O���O���O���O���s`R�Ȼ��Ȼ��Ȼ��Ȼ��Ȼ��Ȼ��Ȼ��Ȼ��Ȼ��Ȼ��s`R�<��O���O���O���O���O���4t��![��                                                ![������t���t���t���t���t���t���s`R�����������������������������������������s`R�R���t���t���t���t���t���D���![��                                                !Z��![��![��![��![��![��![��![��s`R�����������������������������������������s`R�![��![��![��![��![��![��![��!Z��                                                                                s`R���w���������l^�t`R�s`R�l^�����������r�s`R�                                                                                                                s^PIs_Q�tbS�zgY�s`R�s_R�s_R�s`R�yfX�tbS�s_Q�s^PI                                                                                                                        m[Is`R�r_Q�        r_Q�s`R�m[I                                                                                                                                    s`Q�s_Q�        s_Q�s`Q�                                                                                                                                        s_R�s`R�s_Q�s_Q�s`R�s_R�                                                                                                                                        UU+s_R�s`R�s`R�s_R�UU+                                                                    �����   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �� ?�   �� ?�   ����   �����   �����   �����   (       @          �                                                                                                                                                                       [��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![�� [��                                        ![��?z��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��*e��![��                                        ![��k���9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��9v��+f��![��                                        ![��k���:x������������������������������������������������������������������:x��+g��![��                                        ![��l���<y������������������������������������������������������������������<y��,g��![��                                        ![��m���={������������������������������������������������������������������={��,h��![��                                        ![��m���>}��������������������������|x������������������������������������>}��-i��![��                                        ![��m���?����������������������yu������**������������������������������?��-j��![��                                        ![��n���A�������������������yu������%%��������������������������������A���.k��![��                                        ![��o���B���������������yu����������������**��������������������������B���/l��![��                                        ![��o���C�������������������������������21����������������������������C���/m��![��                                        ![��o���D���������������--������������������������+*����������������������D���/m��![��                                        ![��p���F���������������������������������������22������������������������F���0n��![��                                        ![��q���G���������������������������������������������++������������������G���1o��![��                                        ![��q���H�������������������������������������������22��������������������H���1p��![��                                        ![��r���I�������������������������������������������������++��������������I���1q��![��                                        ![��r���K�����������������������������������������������22����������������K���2q��![��                                        ![��s���L�����������������������������������������������������++����������L���3r��![��                                        ![��s���M���������������������������������������������������22������������M���3s��![��                                        ![��t���N�������������������������������������������������������,,����������N���4t��![��                                        ![��t���O�������������������������������������������������������������������O���4t��![��                                        ![��t���O�������������������������������������������������������������������O���4t��![��                                        ![��t���O���������������s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�������������O���4t��![��                                        ![��t���O���O���O���O���s`R���������������������������������s`R�![��O���O���O���4t��![��                                        ![��t���t���t���t���t���s`R���������������������������������s`R�![��t���t���t���D���![��                                         [��![��![��![��![��![��s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�s`R�![��![��![��![��![��!Z��                                                                r^Q&s_R|s_Q�s`R�r`R8r`R8s`R�s_Q�s_R|r^Q&                                                                                                s`Q�s`R�s^Q<s^Q<s`R�s`Q�                                                                                                        s_R�s`R�s`R�s`R�s`R�s_R�                                                                                                        UU+s_R�s`R�s`R�s`Q�UU+                                                                                                                                                                                    �����  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ����������������(      0          `	                                                                                                                               [��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![��![�� [��                        ![��?y��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��$_��![��                        ![��j���8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��8t��*e��![��                        ![��k���:w��������������������������������������������������:w��+g��![��                        ![��l���<z��������������������������������������������������<z��,h��![��                        ![��m���=|����������������������JH��������������������������=|��,i��![��                        ![��m���?������������������)(����EC����������������������?��-j��![��                        ![��n���A���������������)(����ur����¼������������������A���.k��![��                        ![��o���C�����������)(�� ����������##��EC������������������C���/l��![��                        ![��p���E�����������ur��������������������ý��������������E���0m��![��                        ![��p���F�������������������������������##��ED��������������F���0o��![��                        ![��q���H�������������������������������������ÿ����������H���1p��![��                        ![��r���J�����������������������������������##��ED����������J���2q��![��                        ![��s���L�������������������������������������������������L���3r��![��                        ![��s���M���������������������������������������#$��ON������M���3s��![��                        ![��t���O���������������������������������������������������O���4t��![��                        ![��t���O���������������������������������������������������O���4t��![��                        ![��t���O�����������SPP�SPP�SPP�SPP�SPP�SPP�SPP�SPP���������O���4t��![��                        ![������t���t���t���SPP�������������������������SPP�![��t���t���D���![��                        !Z��![��![��![��![��SPP�SPP�RPQ�SPP�SPP�RPQ�SPP�SPP�![��![��![��![�� [��                                            PPP0ROO�SPP�SOO{SOO{SPP�ROO�PPP0                                                                    MMM
SOO�SPP�SPP�SOO�MMM
                                                                            ROOWRPP�RPP�ROOW                                        ��� �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � � ��� ��� (      (          �                               [��![��![��![��![��![��![��![��![��![��![��![��![��![�� [��                    ![��?y��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��)d��![��                    ![��j�����������������������������������������������)d��![��                    ![��j�����������������������������������������������)d��![��                    ![��j�����������������������}y����������������������)d��![��                    ![��k�������������������������������������������+f��![��                    ![��l�����������������yu��21��TR������������������,g��![��                    ![��m�������������yv����������������������������-i��![��                    ![��n���������������������������22��US��������������.k��![��                    ![��o���������������������������������������������/m��![��                    ![��p�������������������������������22��UT����������0o��![��                    ![��r���������������������������������������������1p��![��                    ![��s�����������������������������������22��UT������3r��![��                    ![��t���������������������������������������ZY������4t��![��                    ![��t�����������������������������������������������4t��![��                    ![��t�����������������������������������������������4t��![��                    ![������t���t���t���SPP�SPP�SPP�SPP�SPP�t���t���t���D���![��                    !Z��![��![��![��![����������������������![��![��![��![�� [��                                        SOO�SPP�PPPFROO�SOO�                                                                SOO�SPP�SOO�                                � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 �� ��� (                 @                           [��![��![��![��![��![��![��![��![��![��![�� [��                ![��*f��*f��*f��*f��*f��*f��*f��*f��*f��*f��![��                ![��l�����������������������������������,g��![��                ![��m�����������������������������������,i��![��                ![��n�����������{w����pm��������������.j��![��                ![��o�����������54��������������������/l��![��                ![��p�������������������sp��qn����������0n��![��                ![��q���������������������������������1p��![��                ![��r�����������������������sq��qo������2q��![��                ![��s��������������������������� ������3r��![��                ![��t�����������������������������������4t��![��                ![��t�����������������������������������4t��![��                ![������t���SPP�SPP�SPP�SPP�SPP�SPP�t���4t��![��                !Z��![��![��������������������������![��![��!Z��                            SPP�SPP�QOO�QOO�SPP�SPP�                                            QNNhSPP�SPP�QNNh                        �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �?  
KeyPreview	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShowPixelsPerInch`
TextHeight TPanelPanelLeft;Top Width|Height�AlignalRight
BevelOuterbvNoneConstraints.MinHeight^TabOrder
DesignSize|�  TButtonOkButtonLeftTopWidthlHeightAnchorsakLeftakTopakRight CaptionOKDefault	ModalResultTabOrder OnClickOkButtonClick  TButtonCancelButtonLeftTop(WidthlHeightAnchorsakLeftakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonCheckAllButtonLeftTop� WidthlHeightActionCheckAllActionAnchorsakLeftakTopakRight TabOrder  TButtonUncheckAllButtonLeftTop� WidthlHeightActionUncheckAllActionAnchorsakLeftakTopakRight TabOrder  TButtonCheckButtonLeftTopvWidthlHeightActionCheckActionAnchorsakLeftakTopakRight TabOrder  TButtonUncheckButtonLeftTop� WidthlHeightActionUncheckActionAnchorsakLeftakTopakRight TabOrder  TButton
HelpButtonLeftTopHWidthlHeightAnchorsakLeftakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonCustomCommandsButton2LeftTopaWidthlHeightActionCustomCommandsActionAnchorsakLeftakTopakRight Caption
Ko&mmandonTabOrder	  TButtonReverseButtonLeftTopWidthlHeightActionReverseActionAnchorsakLeftakTopakRight TabOrder  TButtonCalculateSizeButtonLeftTopBWidthlHeightActionCalculateSizeActionAnchorsakLeftakTopakRight TabOrder
  TButton
MoveButtonLeftTop#WidthlHeightAction
MoveActionAnchorsakLeftakTopakRight TabOrder   TIEListViewListViewLeft Top Width;Height�
OnRecreateListViewRecreateAlignalClient
Checkboxes	Constraints.MinWidth� DoubleBuffered	FullDrag	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedParentShowHint	PopupMenuListViewPopupMenuShowHint	TabOrder 	ViewStylevsReportOnChangeListViewChange
OnChangingListViewChangingOnClickListViewClick
NortonLikenlOffColumnsCaptionNamnMaxWidth�MinWidth CaptionLokal katalogMaxWidth�MinWidthWidthd 	AlignmenttaRightJustifyCaptionStorlekMaxWidth�MinWidthWidthF Caption   ÄndradMaxWidth�MinWidthWidthP MaxWidthMinWidthWidth Caption   FjärrkatalogMaxWidth�MinWidthWidthd 	AlignmenttaRightJustifyCaptionStorlekMaxWidth�MinWidthWidthF Caption   ÄndradMaxWidth�MinWidthWidthP  OnAdvancedCustomDrawSubItem!ListViewAdvancedCustomDrawSubItem	OnCompareListViewCompareOnContextPopupListViewContextPopupOnSelectItemListViewSelectItemOnSecondaryColumnHeaderListViewSecondaryColumnHeader  
TStatusBar	StatusBarLeft Top�Width�HeightHint9   Klicka för att markera alla åtgärder av den här typenPanelsStylepsOwnerDrawText'   Fullständiga synkroniseringsåtgärderWidth_ StylepsOwnerDrawTextNya lokala filerWidth_ StylepsOwnerDrawText   Nya fjärrfilerWidth_ StylepsOwnerDrawTextUppdaterade lokala filerWidth_ StylepsOwnerDrawText   Uppdaterade fjärrfilerWidth_ StylepsOwnerDrawText   Gamla fjärrfilerWidth_ StylepsOwnerDrawTextGamla lokala filerWidth_ Width2  ParentShowHintShowHint	OnMouseDownStatusBarMouseDownOnDrawPanelStatusBarDrawPanelOnResizeStatusBarResize  TPngImageListActionImages	PngImages
BackgroundclWindowName2Total actions counter on synchronization checklistPngImage.Data
x  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?0222 ��,F�� ����7���,ׇ̀����@*(�Q�P��oذ6�3c�3�g����71`�:� F�#��٢���79��Ǘ���c5�7I��¡���eH_r�� ��`�.|`K�~$=:�j|�g7�����f�8�1H�c���+�-�f~'�2���bx��v�B��1�p��L�w3�6cx��=v�D���}��9���bb{��{����"����d���a`f�P]�7h���ڔ��ۏ����c��f�9���ɦ����0�fp>x��CT�n�)Ç���`��� �N|���͝� àی���j�O>c7��Ǉ�ߣ��������p��U&�?}�n���7�{/ބt�ژ�������b |��Ӏ1�G��1�?��cK�[�� �w��yhM    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
S  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q@�B�v���������N�B���4n\����Y��. �.th���̑���l���p�tb����ٳ�>����O�,F����8ؖG�^2<�|�Sd 33��˗�=��*���z�P�%1�^�8)�ƁO�n  䳚w�]��    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
X  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q�̑��������*�;�d�B�p<3�4%��W�2<�|�H�RR\l�?�������2�g��pt�I���B���؀=z�a�;[t1F�v�c�
ʖ��:��~c���� ��93q�M�N��*F��� T|��
��@1Kt1���h��8�  �e�dI���    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
R  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q@��Y����32
0������u������@^����g���������B�@��@���H��϶8����0|��̭���~_��Û2�X�_���q��`��`����p��C��O����G��@���;���%1�^�8)�ƁO�n  Ͳ��<�s�    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
R  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q�̙�ã���i��i�?;�d�L^�xff�i:b"\_�bH����(fJIq1|�<���3�XQ������7����{����P�]�蘜�����<�o�?}A6�X�_���Q� �^8
TgR���>[��Q�G����7  �P>�֠    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
v  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�KLSQ��>z���ii�
mx*A�+$l\FcܰacK01х_�.\ibԴcdc4���Mc"�GRT�h�1��}Ж>���� .<�33����?���P*��(��[��~��G��l�|���g2��&J�GNJ҄�3����/܍��ӡ��J�v{Dq`mq?B�<�!�k�A��
����G�\�oF��8+ �$ax$�K�f��HҐZ|���h�
�V;��Z�0��gA�� >tحG[v6 I��(�Hp<���S:]�ٗ;ꪜ��
�����\0�7��..��1Eq1�߳!Ե��X��eA�W�2�������R�/��td0�{%)��W�2 �@�TTt����X��q��ߢ1x?=�����Gԧ�(?�/��W�U���鴻2M0<%�y$i���	 uq}����Z��n&��O?��Ц��)�t�ճ���2�'݅��6��9�"��4�N--�� >��|�\k%;6Wr9x�S�3{l%�|L����$u� ���-躉a��E8�ƴ�������Mڄ�y3"f�8�d���<!����R0�r��h��������(��Wo�����wRp�v�N�R)�f�>�֞_ s'xp�r_�y�0\%�k��3�k �����H��\�8��G�:�,In�W��n�����
%�>%����u�&��������������'�zn�K��    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
v  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�KLSQ��>z���ii�
mx*A�+$l\FcܰacK01х_�.\ibԴcdc4���Mc"�GRT�h�1��}Ж>���� .<�33����?���P*��(��[��~��G��l�|���g2��&J�GNJ҄�3����/܍��ӡ��J�v{Dq`mq?B�<�!�k�A��
����G�\�oF��8+ �$ax$�K�f��HҐZ|���h�
�V;��Z�0��gA�� >tحG[v6 I��(�Hp<���S:]�ٗ;ꪜ��
�����\0�7��..��1Eq1�߳!Ե��X��eA�W�2�������R�/��td0�{%)��W�2 �@�TTt����X��q��ߢ1x?=�����Gԧ�(?�/��W�U���鴻2M0<%�y$i���	 uq}����Z��n&��O?��Ц��)�t�ճ���2�'݅��6��9�"��4�N--�� >��|�\k%;6Wr9x�S�3{l%�|L����$u� ���-躉a��E8�ƴ�������Mڄ�y3"f�8�d���<!����R0�r��h��������(��Wo�����wRp�v�N�R)�f�>�֞_ s'xp�r_�y�0\%�k��3�k �����H��\�8��G�:�,In�W��n�����
%�>%����u�&��������������'�zn�K��    IEND�B`�  Left0Top�Bitmap
      
TPopupMenuListViewPopupMenuLeft�Top� 	TMenuItem	CheckItemActionCheckAction  	TMenuItemUncheckItemActionUncheckAction  	TMenuItemN3Caption-  	TMenuItemCheckAllFilesinThisDirectory1ActionCheckDirectoryAction  	TMenuItem!UncheckAllActionsinThisDirectory1ActionUncheckDirectoryAction  	TMenuItemN1Caption-  	TMenuItemReverseItemActionReverseAction  	TMenuItemMoveItemAction
MoveAction  	TMenuItem
Calculate1ActionCalculateSizeAction  	TMenuItem ActionCustomCommandsAction 	TMenuItem    	TMenuItemBrowseLocalDirectory2ActionBrowseLocalAction  	TMenuItemBrowseLocalDirectory1ActionBrowseRemoteAction  	TMenuItemN2Caption-  	TMenuItemSelectAllItemActionSelectAllAction   TTimerUpdateTimerEnabledIntervaldOnTimerUpdateTimerTimerLeftPTop�  TActionList
ActionListLeft�Top� TActionUncheckActionCaption	Avmarkera	OnExecuteUncheckActionExecute  TActionCheckActionCaptionMarkera	OnExecuteCheckActionExecute  TActionCheckAllActionCaptionMarkera &alla	OnExecuteCheckAllActionExecute  TActionUncheckAllActionCaptionAvmarkera a&lla	OnExecuteUncheckAllActionExecute  TActionSelectAllActionCaption&Markera allaShortCutA@	OnExecuteSelectAllActionExecute  TActionCustomCommandsActionCaptionEgna ko&mmandon	OnExecuteCustomCommandsActionExecute  TActionReverseActionCaption   &Omvänt	OnExecuteReverseActionExecute  TActionCalculateSizeActionCaption	   B&eräkna	OnExecuteCalculateSizeActionExecute  TActionCalculateSizeAllActionShortCutA�  	OnExecuteCalculateSizeAllActionExecute  TAction
MoveActionCaption&FlyttaShortCutu	OnExecuteMoveActionExecute  TActionCheckDirectoryActionCaption(   Markera alla åtgärder i &denna katalog	OnExecuteCheckDirectoryActionExecute  TActionUncheckDirectoryActionCaption*   Avmarkera alla åtgärder i denna &katalog	OnExecuteUncheckDirectoryActionExecute  TActionBrowseLocalActionCaption   Bläddra &lokal katalog	OnExecuteBrowseLocalActionExecute  TActionBrowseRemoteActionCaption   Bläddra &fjärrkatalog	OnExecuteBrowseRemoteActionExecute   TPngImageListActionImages120HeightWidth	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  BIDATxڕ�KLQ��J�U4��S. E�"�T���
���Ԥ	�Pe�N��+���$$���mm-DcecX��MD1X�}"	��v"#M;��_�9s�wO�d(�a����+C�-��LZ�\O�r�l:T>�`H���1̶I�5H�.Q��y�%(�mm49>e2�Agb`^_q��`��;;���r��CY��[�{;����郩�`ӹv�S߁�LX�!�-"�m�-��.��6�K/|XB���p���<ۆR�	I��B��*��d�U~���i�����.��Fq�Ax�G	G���6v���N�L)G�N9<<�j�X��'N�b�&7�eb��F4y�QTQ�ּ}Ո���AU���76�BRW�M�Uՠ@*C퐓���b�?��� �ؐ���Mf������fM��������#`<� �Z�h�ϟG����Y��>�Ki����F"��jv����j��f~�T �[�c'�T!�Z�k��(��36}}:�����g}(�!��\�uv�M�",�{�b2�[%�)+C,�]4�� (�R�il�7&G�xz��)R��쌣    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?5㨁�H��v�������������u�Th�����p�������|T�a!�:{82�����¹�_�|Y��绬g��ʷfd`��i�����������a�2�20�+W>z|��ϯ`P0�ș��]���K������defe`�O�<e8s����$S�@�ŋ����D}��(0�����P�%.q�aH�X�Pp?P� Μ2��Ao  �?�ƻ�1�    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  'IDATx�c���?5㨁��MP�IH������/T����@�6�x�����.]gxP���,���؅������3�s�1�ݱ�<�y4X�����j��h3����~�Th:	Ti��=+߹bgTh�dbf�kb`�)-#��h�￿Ql�/g&wţS/q��?�Y��IH�����Tv!,Y����ɪ����?jʷ�cd`4D
�}�0t�&�A�.v��||���zl��22�oJfae�
L��W/^��@�i�cabX��w�$8��Ao  �S�
G�j}    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?5㨁�H���<{���c�����:�����o '�p��������L��u!��j3|���̝���X���sV:�7��3yy302��u��$��[��PYY�213\~�����W���g#H�\߮_��?}�+3���X��~�p�����I��� ����N����.��=
�+DP1������8�0�z,x:��˳�?#� Μ2��Ao  r^䭱"�B    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?5㨁��Mp*�&�2�]�2>q�������L�L��d�9/<zʐ��3#Y�d`�b�����o������̰��U�{��a�����������8���0#�\��c�?[cg������2�@S�SFT����?@�P������׷��/�� ���ƺ`C(6��.$.y�UZ���?É�ϟ-���&�i��,� �����_lI2p���@ ڎ�f+��    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
P  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڭ�[lU ��̙�vn[6K���K)�*.�n@c$$_������`���}0��XJ5�Ã�}2*��DYV@H�B��.t�nwq����g<3++�T|�<����wr��̏<σ�9�"������$�^R���Y���$)� �l+�W� J`�}l�,�����[�({i�\���[�ç��-��B�&d߀�)�B��;�ۻ.^��L&�}���(�ދKR�C��D"mm{R�������	�Ѱt(R�rw�.�,�u��K��������F��|�p?v&�ubp��\HO�2�kHU�pD��
�8ٹc��P>tR-�.}|XQ�
������s�v1��b� ��Sy�u�R��9�����M��� �m���P$������p_w?�����p�H 51�����@I;�_�cD�iǈ�9����h� fZ6����u���$<��ɉi˰�T��t���c��7lkojb�Y)6
A�0!9u��-�@����]���*���O��H�>�ϼaY��:e�z�B>���k�����"B�+�-M�&�5~��1�~n�h��R,D��b"�b����rk��<�߹�Ţ�zO���O�(��������Iz-��?>����(�]�h:��9��կ��+y��[a���T��K�U�����U�~��n�Q4C���Ҝ�x݃�����ƿlj�7B���
C?�-)����n�.�����2�b�5���I�({�(T��dy(±�t��bWu�����~'�vY~���S�D�]�Y�Z�F�����Xܷ����mÌeф�g����H�����YG���a@�q����j+���3�o�s�L��=R.ϯ�Eq_3cM#�9Nζ�~M����X�M�>���݄�c<�Ű��Ę���a��(���祂e    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
P  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڭ�[lU ��̙�vn[6K���K)�*.�n@c$$_������`���}0��XJ5�Ã�}2*��DYV@H�B��.t�nwq����g<3++�T|�<����wr��̏<σ�9�"������$�^R���Y���$)� �l+�W� J`�}l�,�����[�({i�\���[�ç��-��B�&d߀�)�B��;�ۻ.^��L&�}���(�ދKR�C��D"mm{R�������	�Ѱt(R�rw�.�,�u��K��������F��|�p?v&�ubp��\HO�2�kHU�pD��
�8ٹc��P>tR-�.}|XQ�
������s�v1��b� ��Sy�u�R��9�����M��� �m���P$������p_w?�����p�H 51�����@I;�_�cD�iǈ�9����h� fZ6����u���$<��ɉi˰�T��t���c��7lkojb�Y)6
A�0!9u��-�@����]���*���O��H�>�ϼaY��:e�z�B>���k�����"B�+�-M�&�5~��1�~n�h��R,D��b"�b����rk��<�߹�Ţ�zO���O�(��������Iz-��?>����(�]�h:��9��կ��+y��[a���T��K�U�����U�~��n�Q4C���Ҝ�x݃�����ƿlj�7B���
C?�-)����n�.�����2�b�5���I�({�(T��dy(±�t��bWu�����~'�vY~���S�D�]�Y�Z�F�����Xܷ����mÌeф�g����H�����YG���a@�q����j+���3�o�s�L��=R.ϯ�Eq_3cM#�9Nζ�~M����X�M�>���݄�c<�Ű��Ę���a��(���祂e    IEND�B`�  Left� Top�Bitmap
      TPngImageListActionImages144HeightWidth	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   IDATxڵ�ILa�w8x1F��A5���a�%
����`P�����xr�q�J���Ph(�qI4XhK�R��@�;N��b|{����=g�EQXA�O�M/�u�ӗ���Ty�u�������[g���. �t�X,��3����(�/�^;O�^���m�����D�U�'C�@ ������A�b��1�v��>��TF��Pܼ<L�Y�jEJ���\�֕��p����=�R�)PP�Ox��FuB�k]���L0����u��cH��~ظ:��W_"{)� s����*ؓ_ y�*��,C� �E��SSda�>	oj �Rj`К���L�?A�f�*��v�I���z��>��0�xN�C7����q�����DpF^~�A-�:33����H7ȳb���WB�_-AB�["���3.�U#0�-��Z���<�^����E����)Z�f���O�a��d���d�J�s
�v�z�_!�V��Z	v���B���l����{�+�B#33h�
���o����&v�w� �����@�5�b�y�P������MhThK�`n�YP�#���#���ã0�a��2��4��;A^j^�;������n��?H�Ao��:�Ĥ�a�K
���m��F���B�--�F�ϵ�����m����\
��V�ٽD�[0:��NM�@�w�J>��I��b�ؘ��JI�R�����X�6��'��mAA��uk���zvv�	�L��k���KA�������}���O�    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
-  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���KQ���B��K7���B�����d;�%<F@At��:T�c5��Q�vX�窻�+�N����B�D���=���y0ߙGFi�����&v�Cn&�ғ� �Q���y<U�z �8Eq0�����< e$-\�Ᵽ���"�]�h	���i�~�N7�-@0:qF�̵'#�)���� Z �����u�UN��F``z��uҍB������d9�8�t}���q��>[��-�[�rd�X"RN�vPȿ���0�=��H��v!g�Dre_2��� $�J�A�K��EvB��b��ɦL+u�E9(�d:��h�v��v������V����^�wLU�C���2�7̰[&�bz��������u�"Yi��/    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  lIDATx�c���?-�o!r��� �Q���T�@�A@�?;�$nn��o_��zP���j�\���<O^^VFIU�����*��-A��X�;999s��u�����ðw��-Ph���ļD^^NY[[��������?(ȷ�jpA3�P��#C��`#{���	���ß��-Ph�/g&�b£S/��%��J�9��00�03�Jm�J�ۙ�Ȃ��l��������"G�M�������pE�^�'dC�3�?���.9�d�&4���3YO_�����ȶ
�331,�S�WVSdؿ�u- hQ1���;�ۗ��-*��|�����.�~}0j!  �\�?'(    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
&  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  }IDATx���KA��Т���DעNQ�蟐@�Qޢ?"�塿 :t��t��NZh����mAsg�]W�i2WD�V"�]��7����7�c�KC}���-��zg�քeJ�{�Tt��H��_Ԉ��a����F�AV!��JY��x�(`a|�_� ���P�ثb��
@ꀐ$�BS�j���L��5 � @��b�4���	��b���o O�s�lk��&4�1���J� 7wq���m�-���2o�H�2Y��g���8�3ʵ� ��A8�Č���%d��,]�^���WKO��5�A4��%r��쫋�D������651�h��Am�>h��X��d��y�$Q�=� �*�7�ݬ5��Vσ����>��}�f~N"    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data

  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  aIDATx�c���?-�o!3��]At�ׯ��jA?� /�$��/?~�J����j�\���8OA\DFSB�aۥ��>�-Af20p1��tr���(�3ss20��˰��U�-���i����DNBTY[A��(���f�� ��� `9����%.9�6I^�Fv6�r-UFqA�����wccCq�_���1����/))栯�����4�/u-���sPJR̎f ��C�������P_K��A�d^^[fF���HV�ɠ����耚N��O����F2���=���#�PI�A���L��vgfb\�h�T�h� TTp��L�eg��zQ���qy2�e�Cva7��Q (� �?�Y�    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  ;IDATxڽ�{lSu��������Q�X"8P���GV���?��Pb�1$&v��@�CL��`|�W2Ɔ,F_!�DM �âs�B��	��l����{��{{{=�k���<Iӛ_�9�s���;Ķm��F�7 !d��[��4Н`��Z�׵&: �M��~	+j�;��) d�8�=�u�fall\�LkG���[-y��|��������]�����@\i]薝M����PV�p8C��Eӆ�E�/����,��`��F[R�H$
�����%�C.9�P�uo(_�M�a$x!�c'��Ta�b_T�y���H� ��A���i�VU=� K=�b����!`&�d|r
��|]�;�͝���ے��l�������غn>ע�?�G���$��G�>�~�Z/p,���^������(;o $�E�3�$t4�<8���Z��)ʗ٘@NE�������7UW���/N��L��+�v�/�� M�`���[p-�&v�A�E�B��<�v��m!���E��	�2h��E��,���}ڪ(�-����!��<�1_��lbKDai�f�O#02��a�/�*�U9}3�}��
�#����l�L��\W�g�������9Y�)ݴy�;���LL��oa��/�>Vt���%p̻~]��b� ��F��i�L+��5�������=����ڕ9W����ɬ����)+��MU�	����a�#��b��;��Z��B�_�O�U]��	3��ae�l״��gX�|�PR�s�=���#���^b8.�GG+������a؜��fs{<9�,��,����s�Dd�|�Xᙸ���֣m��H�� ����e�D�0[����ըnۏ����.Y�9y�d���ZN������W���4�rY���fv��c��b��de�$�[ R��P_�p=8�Y�{:���y�%��y9)"���㢨��1�Ÿ�x�s����;葄�<�>��.��i����k_�*�+��E��W�q!�z"�
���˪(��Q)��\�]�%��:�#�"fk�fW|wj�Ge$����K\�ݲ �1�'-&    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  ;IDATxڽ�{lSu��������Q�X"8P���GV���?��Pb�1$&v��@�CL��`|�W2Ɔ,F_!�DM �âs�B��	��l����{��{{{=�k���<Iӛ_�9�s���;Ķm��F�7 !d��[��4Н`��Z�׵&: �M��~	+j�;��) d�8�=�u�fall\�LkG���[-y��|��������]�����@\i]薝M����PV�p8C��Eӆ�E�/����,��`��F[R�H$
�����%�C.9�P�uo(_�M�a$x!�c'��Ta�b_T�y���H� ��A���i�VU=� K=�b����!`&�d|r
��|]�;�͝���ے��l�������غn>ע�?�G���$��G�>�~�Z/p,���^������(;o $�E�3�$t4�<8���Z��)ʗ٘@NE�������7UW���/N��L��+�v�/�� M�`���[p-�&v�A�E�B��<�v��m!���E��	�2h��E��,���}ڪ(�-����!��<�1_��lbKDai�f�O#02��a�/�*�U9}3�}��
�#����l�L��\W�g�������9Y�)ݴy�;���LL��oa��/�>Vt���%p̻~]��b� ��F��i�L+��5�������=����ڕ9W����ɬ����)+��MU�	����a�#��b��;��Z��B�_�O�U]��	3��ae�l״��gX�|�PR�s�=���#���^b8.�GG+������a؜��fs{<9�,��,����s�Dd�|�Xᙸ���֣m��H�� ����e�D�0[����ըnۏ����.Y�9y�d���ZN������W���4�rY���fv��c��b��de�$�[ R��P_�p=8�Y�{:���y�%��y9)"���㢨��1�Ÿ�x�s����;葄�<�>��.��i����k_�*�+��E��W�q!�z"�
���˪(��Q)��\�]�%��:�#�"fk�fW|wj�Ge$����K\�ݲ �1�'-&    IEND�B`�  Left� Top�Bitmap
      TPngImageListActionImages192Height Width 	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx���klSe����Ic�(š��,xL6�A��k���m�B�ױ1����ۚ���Eg4�l�m�q��F�1�u��{z[/(^�oO�����R��S�^���?'M��B�?�����^z��x�����CI�;��.8[;z�����%�u3 yyu�;�;�wix� d�frbQ�
r����O�X�>m��?�ʪ!{[ȍZr��2��A��Ork/��u�g��� -�gx�=�������R��љ`:�_L�r��.����^�B�jO���=,������0�PvL�=ڤ �Y���ه�V�2)��V�xβ��`cu� s[Wt�E�W�e{}��H�,5�2E'R����� ­�4�S 8M:��4�ZY8����ii�=Oe��I=`�9�F�o�O'�zVe�7�Gn�'�ɠm��4e������^�`;w����[+�p1�sj��Ҡ=$�y�
����Xf� �ݜ���`�g5��Pi9��m-�y�
��C�{N����4��ۍ3�H���H���Yx)���O��^N鏯���
KKʣ[�1�F;�-@.�mr��o0���H���?Gӳ��İ�p;)�ȋ`����?�f%�$��*d���lk>,����5GX+������o�5f�G�wW"sﻸW�!z��wg�W`�|����}7�aa�q�(R	,:-�E 3_u@���KOǊCG"�Mjm6�=��o/����~@ 6'���5E�/j |�xt}��Z�[��,��r�2��x��_�@|z�4o cwa�C��4����D��AL\E̿�n�f�!��	K�g��*Nx�t�Յb�.��`�ɸ��wja �p����'N��Dp2n��t�\0��@Xu2a��}0|܌�ͭX$��_5M���=��hb1f��V��n��-��JӰn�~�PP��0��G*�=�����(9�6aZ��5�Sh�����!�DX��S~��^�AJ�}K��1�-�+x�W@� �Zy˦�RvLes����K��F�1�    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
e  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���MKA �w���nյ�SP]�Eu��QVx3:��~@t�����4
uM�]Bpu�Rv��f#��C�^v`�a���g�yw1��Ά�p ��:ag�{��a3�ϸ��
xYo7$bul�5�*n��T���Xfb�q����I���I���wd�'P�J2�Y6v�:�h�Y2�T[*��y�q�n�]nx}�B8�R���L:��� t�7}�L0�R5�� F��h,��T�R2����(���y��Y�Z���( �PEB�f�[ �2���@:����u��k�֪�R�@¸��C2��;0����!/�3~s��K�xHLZ���#��{�ĳO�r��P΋HIT(�겱�5�� uC�.��N?L'��R�Y�� �z@�&��׬�䏑�gm#��eWJ�����!q ��x��|O3�Z�    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
`  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?�@�Q�:`�� bɶ
�033,��������s@��@3+K�����7T�#��;@�EH���a�������;+���� �v�H&&��jj�
J����⿴w�B���v�i|���FFF<����e�����B��l��g��V��Qw�\+�3#3�U%e--M��b\Ph�/g&��W�N�$Z#0��)pu����[�3����-�YLs ���������)33�2�:@� ��r@�P;G������� %21/VUV���Ҡc"D�l���4���7��А�O6F�~`.v�f0�v9���	1�*rm�,��S�5�y�d�W!�y6&���"B�Z�t.�� Xɳ	��2�ih��^�x����VA=f���`FUx�d��u�@;  9�P[��    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
n  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�햽K#AƟɊUV�Z��F�:���?AAIDE��$�Xj�6� �*"r~���qzhL��Lfg���θ�;4b�s��if�y�1�;�;D?	 � �w��m8���	A�툞���LU����)�r!F�)�\*@GcL��^�
w�jYv��i&�@	��B����IB��;C�f� L�� ����k�������(�@��}z��n�T��
<�p�WV��],�R�b\��5 �P ��<��Oji�EW��%� (�C��b��T�r��k]�.�۳����4-�������?Hi7?� C� g��RC�%��e
�	-�p�����s��[ZJ�7���KѸ\ݻ����{����rVJ!��Ԩ�8�Q�f^�? ��^z�X�(XV�i�K�?�����b3���h4&�M��AP-l�5�_���� @ �7�F��32.    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
f  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��AKQ���[w�}OSH]��"�42�]�Ry�}��D��]=�`%TT�:Dt�+D?Ab�
S_O#)4�����mav��f���C�0  �� �$�	�Ny��{-�%�
��Ȏ���y��s�}��[��K�Қ��.���2DVYF�OY1 ǔ�I:�1���sR�t ��M��P��7gB#�n���J�	��� ���=�
�X����k ��e^���u"��#�X��'@������h�TB�U�QpJE�d_UL{�H�NG�X��������x4D
ƍbȝ��Z�
�8�$�ځYUw�
�݂�#B������k�"V�F���f��o����Z!���ك܈�(#�5+6a��Ӵ�o�E�bj�%�t�� %#>]�1��?����s\�M��9���`  ��uӻZ��h    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
6  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��[lSu���sz;�t���:W�F.[W��Q2�����KI���<�4�| AtL�����@@�1`���Vƺ[��������e��݌�/M�������~��A�,��4��@�k�v������ߜ � �b�dT���.�y+��B*x?!�4���s$������F�� ���6?�����B?8Ǹ�ڵ�/tBp�����;r�7���j�� Tp��*ܾ�?�!^���<���X�Pq�eC�k%$�pN�:����]Y�
Кt���ν:�)�����/p�n������ i`~(-�ֻV9�T 'p����G�j����F`B���<�F,Cg�pC�������Y�.��8�Ȓb�J�C��r�������� ��r���2�6�V������$�Y1��5��3��t6 ��
�s�c����kA��)�|]J�Y���@��%�o�\��2�N�x�^�P(����}��/XM%���N{y��V�^�����m"ǽ��OGt�2l5�בu�f�Cg1�e@D�18��CB�-���V��
g��K+�eVKz���7�����<Ȑt.�d2��:��:Q娠�ͦ�9g���?�(�$Th���N[�����a���b��)�.׼ ��0N
��V�m�2�9cn�C�Tc�͆R��K7n�H�1��-Y���C����:����VQdɘ�pu��R�����%D�)O(�9lA ����hH�g{a�sY�5�	,�_$*	k�r�6�����q���a�=^�)�(%�̍���w �4�]d`>3j���PČ5���׆��f�?hV�����@�{Յ�?U���g`zG'�%�{~j�/ ��Y���֭�*,�X�$�wd���D�j`8>��-
`�Qϲ�J}�
�Ƨ��fC��E�j,��|���߅����?ǿܜ���O�_�}`���p����zߋƾ�O�[E,���$?u�����\��h�@ڼ ��Bgc����w��A#1��`=����g�M�:P�oB,uBR ��q���8)��@�|jg�mY�����z(������O׷�e7P ��3P&�J��q�\���(m��g�!=���*Zg�N0�|��F�E�:W���z�P��R��-�g���HBN��� "�.f��J��Y���p]zA�ڹj�E�s�$yܩ՘K&�`��pX�&�-<$�-S�Bp�AQ����~Q�A���]�'�yX�S�OK)��6��<�h��b1�/l��`�$LC����c]qq$&��n�y�|����y�N�v�'��w$Iɟ5;eY�	0B�Pyĵ��H�B��!�rF�/RU�	9�e4�FԌ[p! �0��)S�)a�ף`� ��ex�?���3����H    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
6  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx��[lSu���sz;�t���:W�F.[W��Q2�����KI���<�4�| AtL�����@@�1`���Vƺ[��������e��݌�/M�������~��A�,��4��@�k�v������ߜ � �b�dT���.�y+��B*x?!�4���s$������F�� ���6?�����B?8Ǹ�ڵ�/tBp�����;r�7���j�� Tp��*ܾ�?�!^���<���X�Pq�eC�k%$�pN�:����]Y�
Кt���ν:�)�����/p�n������ i`~(-�ֻV9�T 'p����G�j����F`B���<�F,Cg�pC�������Y�.��8�Ȓb�J�C��r�������� ��r���2�6�V������$�Y1��5��3��t6 ��
�s�c����kA��)�|]J�Y���@��%�o�\��2�N�x�^�P(����}��/XM%���N{y��V�^�����m"ǽ��OGt�2l5�בu�f�Cg1�e@D�18��CB�-���V��
g��K+�eVKz���7�����<Ȑt.�d2��:��:Q娠�ͦ�9g���?�(�$Th���N[�����a���b��)�.׼ ��0N
��V�m�2�9cn�C�Tc�͆R��K7n�H�1��-Y���C����:����VQdɘ�pu��R�����%D�)O(�9lA ����hH�g{a�sY�5�	,�_$*	k�r�6�����q���a�=^�)�(%�̍���w �4�]d`>3j���PČ5���׆��f�?hV�����@�{Յ�?U���g`zG'�%�{~j�/ ��Y���֭�*,�X�$�wd���D�j`8>��-
`�Qϲ�J}�
�Ƨ��fC��E�j,��|���߅����?ǿܜ���O�_�}`���p����zߋƾ�O�[E,���$?u�����\��h�@ڼ ��Bgc����w��A#1��`=����g�M�:P�oB,uBR ��q���8)��@�|jg�mY�����z(������O׷�e7P ��3P&�J��q�\���(m��g�!=���*Zg�N0�|��F�E�:W���z�P��R��-�g���HBN��� "�.f��J��Y���p]zA�ڹj�E�s�$yܩ՘K&�`��pX�&�-<$�-S�Bp�AQ����~Q�A���]�'�yX�S�OK)��6��<�h��b1�/l��`�$LC����c]qq$&��n�y�|����y�N�v�'��w$Iɟ5;eY�	0B�Pyĵ��H�B��!�rF�/RU�	9�e4�FԌ[p! �0��)S�)a�ף`� ��ex�?���3����H    IEND�B`�  Left8Top�Bitmap
       TPF0TSynchronizeDialogSynchronizeDialogLeftoTop� HelpType	htKeywordHelpKeywordui_keepuptodateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"Keep remote directory up to date XClientHeight�ClientWidth�Color	clBtnFace
ParentFont	
KeyPreview	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize�w  TLabelLocalDirectoryLabelLeft1TopWidth� HeightAnchorsakLeftakTopakRight Caption.   Be&vaka förändringar i den lokala katalogen:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft1TopDWidthHeightAnchorsakLeftakTopakRight Caption6   ... och inför dessa &automatiskt på fjärrkatalogen:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  THistoryComboBoxRemoteDirectoryEditLeft1TopTWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeft1Top#Width8HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeftoTop!WidthKHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButton
StopButtonLeft� Top8WidthXHeightAnchorsakTopakRight Caption&StoppTabOrderOnClickStopButtonClick  TButtonCancelButtonLeftTop8WidthXHeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  	TGroupBoxOptionsGroupLeftTop� Width�HeightwAnchorsakLeftakTopakRight Caption   Alternativ för synkroniseringTabOrder
DesignSize�w  	TCheckBoxSynchronizeDeleteCheckLeftTopWidth� HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTop\Width� HeightCaption*   Använd &samma inställningar nästa gångTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionBara &existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeRecursiveCheckLeftTop,Width� HeightCaption&Uppdatera underkatalogerTabOrderOnClickControlChange  TGrayedCheckBoxSynchronizeSynchronizeCheckLeft� TopDWidth� HeightAllowGrayed	AnchorsakLeftakTopakRight CaptionSynkronisera vid s&tartTabOrderOnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top,Width� HeightCaption&Bara markerade filerTabOrderOnClickControlChange  	TCheckBoxContinueOnErrorCheckLeftTopDWidth� HeightCaption   Fortsätt vid &felTabOrderOnClickControlChange   TButtonStartButtonLeft� Top8WidthXHeightAnchorsakTopakRight Caption&StartDefault	TabOrderOnClickStartButtonClickOnDropDownClickStartButtonDropDownClick  TButtonMinimizeButtonLeftTop8WidthXHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClickOnDropDownClickMinimizeButtonDropDownClick  TButtonTransferSettingsButtonLeftTop8Width� HeightCaption   Över&föringsinställningarTabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxCopyParamGroupLeftTop� Width�Height2AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamGroupClick   TButton
HelpButtonLeftsTop8WidthXHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelLogPanelLeft TopYWidth�HeightdAlignalBottom
BevelOuterbvNoneTabOrder	
DesignSize�d  	TListViewLogViewLeftTopWidth�HeightZAnchorsakLeftakTopakRightakBottom ColumnsWidth�	WidthType�  Width�	WidthType�   DoubleBuffered	ReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReportOnCustomDrawItemLogViewCustomDrawItem
OnDblClickLogViewDblClick
OnDeletionLogViewDeletion	OnKeyDownLogViewKeyDown   
TPopupMenuMinimizeMenuLeftxTopx 	TMenuItem	Minimize1Caption	&MinimeraDefault	OnClickMinimize1Click  	TMenuItemMinimizetoTray1Caption   Minimera till system&fältetOnClickMinimizetoTray1Click   
TPopupMenu	StartMenuLeft Topx 	TMenuItemStart1Caption&StartDefault	OnClickStartButtonClick  	TMenuItemStartInNewWindowItemCaption   Starta i &nytt fönsterOnClickStartInNewWindowItemClick       TPF0TSynchronizeProgressFormSynchronizeProgressFormLeftOTopBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynchronization XClientHeight� ClientWidth�ColorclWindow
ParentFont	OldCreateOrderPositionpoOwnerFormCenter
DesignSize��  PixelsPerInch`
TextHeight TLabelTimeLeftLabelLeft� Top1WidthOHeightAutoSizeCaption00:00:00ShowAccelChar  TLabelTimeLeftLabelLabelLeft1Top1Width-HeightCaption	Tid kvar:ShowAccelChar  TLabelLabel1Left1Top	WidthHeightCaptionLokal:ShowAccelChar  TLabelLabel2Left1TopWidth)HeightCaption   Fjärr:ShowAccelChar  
TPathLabelRemoteDirectoryLabelLeft� TopWidthHeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  
TPathLabelLocalDirectoryLabelLeft� Top	WidthHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelStartTimeLabelLeft� Top1WidthQHeightAutoSizeCaption00:00:00ShowAccelChar  TLabelStartTimeLabelLabelLeft1Top1Width3HeightCaptionStartad:ShowAccelChar  TLabelLabel3Left1TopEWidthBHeightCaption   Förfluten tid:ShowAccelChar  TLabelTimeElapsedLabelLeft� TopEWidthOHeightAutoSizeCaption00:00:00ShowAccelChar  	TPaintBoxAnimationPaintBoxLeftTopWidth Height   TPanelToolbarPanelLeft1TopsWidth� HeightAnchorsakLeftakBottom 
BevelOuterbvNoneParentColor	TabOrder  TTBXDockDockLeft Top Width� Height	AllowDragColorclWindow TTBXToolbarToolbarLeft Top DockModedmCannotFloatOrChangeDocksDockPos�DragHandleStyledhNoneImages	ImageListParentShowHintProcessShortCuts	ShowHint	TabOrder ColorclWindow TTBXItem
CancelItemCaptionAvbryt
ImageIndex ShortCutOnClickCancelItemClick  TTBXItemMinimizeItemCaption	&Minimera
ImageIndexShortCutM�  OnClickMinimizeItemClick     TPanelComponentsPanelLeft Top� Width�HeightBAlignalBottom
BevelEdgesbeTop 	BevelKindbkFlat
BevelOuterbvNoneTabOrder  TProgressBarOperationProgressLeft1TopXWidthmHeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder  TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeft�Top�   TPngImageList	ImageList	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
u  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ��JA���.��v�R��E!�+d/��
�]hu�+T��EY7]iu�T�P bAY�nQ�;әugYM��\,;3��۝���9tSD !p�iDe���d�� �+�1��]���D�4˶W<u= �C����+c'%�\���Y;R����
���)�(K�eHU"3�b;n" Ҽ��@q\�,(6�+,I@&�дx!�5�k���ƪ�!Dӵ�aJ���-
E�Ͻ1v�7�x��b���k�!B�a4`P �#�󶙟��r��( �$���:p��h�p���L��6@�� Ҭ�y
��i��ၸ �6kh��� �}�t [��f}���㔺�g���CV p-�am?U�m��OI�h^P�Ź�*��c�#Äw��$�(���?(�v̢U���!��2�z��eB�)��8X3פY��T|Z�0�Ŀ��\�n�mB���,    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   %IDATx�c���?%�qԀQ�����xM�g��t �47� OWL    IEND�B`�  Left(Top� Bitmap
      TPngImageListImageList120HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڭ�[K�@�l�]�-H+��"���`�C�L�'��"�~�}�/�"�eETD�n����&�g�,�$��K6�s~�ٙ94�"�
�RښXw�/�g������l�������mɹ���NaѢ�r��0��U��Ұ�Ba�0�����piޫ�$@����#����Jl������  �m�����5�g�Y��ކaU��h����Z���Jm�	n�����O5PGŽ�=��|�[�Vn�,�>��p��;뙬"�(C��$"�y��~kIT�Of��V u�;�Ģ��*:
�KC� ;J�^� ���� ��Jl8g�%�z�_.Y`��!`�
V�E�;J�Eb�%�CbY$bd>ӷ���6v	mJ����2N �;���nlq�,�"�n��5�_i%�*z���8.@|��=���G�o4L]4�~ �p,Л�ھL��/�B�h�g�/9D��������3cղ�r���6���q�� �    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR         ��   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   -IDATx�c���?5㨁��8j�����H�@���5��^t �C�����    IEND�B`�  Left� Top� Bitmap
      TPngImageListImageList144HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڽ��/�@�gZ�Ŷ��AB�F��"qw�pę�
w���_��]D"$B���b���ߩVf�3��Ի�����g��}Cc$Ϡ�&����U��#��2��ݗ��@���:%t�0���y5��ኂN���i:u����y��p���6�J�o|��Y.Ivl;��mk#>�G����>�z�K�_G�E׭5	�%k�l�sc(�#M"������_jx�`���A%��jY��Zb2!��Y5|!�M�W���p ݽ��+�Q2i�	9w��M�LA,)A2!I���S��� SKlHH�~��3�]�kܒ`\#8����-JVFpQr	��Hk��Ë��H� ��sW��H��״��1~��{$JAR n# �ΪQ����� �2h�ƻ  o���B: ���|��Rc�M�s�Gûb���ԋ����G$�]<�!pJh��\��G��!P�k�����@�#.J
���'�#3��]�#����    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   /IDATx���  �@�_�XȖV@�$�2� ��x~^��N�S�{���    IEND�B`�  Left� Top� Bitmap
      TPngImageListImageList192Height Width 	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
p  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���AkA����d���J����A�b+�ă'Q<�$��C꿰�
�Q�^s�x.��VDPPJբb�M6U�3��mv²�ٝ�:��fw�'�Lv��������@).��	%�R�����A&^.�/½"I�k�u���]�4@4��\ղ�z�]!��"0nS�lڶK���m!� b�������l;���"T|⣌���U�w������yW�q�q.}��j��k���������M`����������*9��5K���B�0��$���j=7��=/��.�b���� ��/�Ec��L�^�a����@TR&n�����5����5��(�փ �����DoA��[O��gm;�60�:vŇ�S�(� Zù�	����#�d 0��A�w�Ѐ{�s��N�� � x��>�E�
 ��[�e������g ��I��r�j�0�b ��OB���D����HAT��߀���'a]��L � � ~�#)������{��z�k?BD�\ <���1ƴ�O��q��q�"�ei���9lO@�f�q<���6�/�v+��#� j[B<��@R�d~�z|Ab��&�DM ���#:��Hԑsc�7N�O"�q ����{q�#Y�P:| }7�'����(�dr(M;��o���B������z�������F~ŏ    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
�
  �PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   8IDATx���  1޿�	�Hz����Y           F�\Q�W � �����o��pf    IEND�B`�  Left8Top� Bitmap
              @   4        �      @4   V S _ V E R S I O N _ I N F O     ���   M                                     �   S t r i n g F i l e I n f o   z   0 4 1 D f d e 9   >   C o m p a n y N a m e     M a r t i n   P r i k r y l     n #  F i l e D e s c r i p t i o n     S w e d i s h   t r a n s l a t i o n   o f   W i n S C P   ( S V )     *   F i l e V e r s i o n     1 . 7 7     � 0  L e g a l C o p y r i g h t   �   2 0 0 3  2 0 2 0   A n d r e a s   P e t t e r s s o n   o c h   R e n �   F i c h t e r   < 
  O r i g i n a l F i l e n a m e   W i n S C P . s v   6 	  P r o d u c t V e r s i o n   5 . 1 9 . 6 . 0     8   W W W     h t t p s : / / w i n s c p . n e t /   (   L a n g N a m e   S w e d i s h   .   P r o d u c t N a m e     W i n S C P     D    V a r F i l e I n f o     $    T r a n s l a t i o n     ��                